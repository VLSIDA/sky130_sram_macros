**************************************************
* OpenRAM generated memory.
* Words: 256
* Data bits: 32
* Banks: 1
* Column mux: 4:1
* Trimmed: False
* LVS: False
**************************************************

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_7
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_7

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=6 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=6 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_10
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 26
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=6 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=6 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_10

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=2 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=2 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_9
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 9
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=2 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=2 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_9

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=2 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_8
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 3
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=2 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_8

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=17 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=17 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_11
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 77
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=17 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=17 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_11

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pdriver_2
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 3, 9, 26, 77]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_7
Xbuf_inv2
+ Zb1_int Zb2_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_7
Xbuf_inv3
+ Zb2_int Zb3_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_8
Xbuf_inv4
+ Zb3_int Zb4_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_9
Xbuf_inv5
+ Zb4_int Zb5_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_10
Xbuf_inv6
+ Zb5_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_11
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pdriver_2

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pnand2_1
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpnand2_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_nmos1 Z B net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand2_nmos2 net1 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pnand2_1

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_20
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_20

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_delay_chain
+ in out vdd gnd
* INPUT : in 
* OUTPUT: out 
* POWER : vdd 
* GROUND: gnd 
* fanouts: [4, 4, 4, 4, 4, 4, 4, 4, 4]
Xdinv0
+ in dout_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_0_0
+ dout_1 n_0_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_0_1
+ dout_1 n_0_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_0_2
+ dout_1 n_0_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_0_3
+ dout_1 n_0_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdinv1
+ dout_1 dout_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_1_0
+ dout_2 n_1_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_1_1
+ dout_2 n_1_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_1_2
+ dout_2 n_1_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_1_3
+ dout_2 n_1_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdinv2
+ dout_2 dout_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_2_0
+ dout_3 n_2_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_2_1
+ dout_3 n_2_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_2_2
+ dout_3 n_2_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_2_3
+ dout_3 n_2_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdinv3
+ dout_3 dout_4 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_3_0
+ dout_4 n_3_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_3_1
+ dout_4 n_3_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_3_2
+ dout_4 n_3_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_3_3
+ dout_4 n_3_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdinv4
+ dout_4 dout_5 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_4_0
+ dout_5 n_4_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_4_1
+ dout_5 n_4_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_4_2
+ dout_5 n_4_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_4_3
+ dout_5 n_4_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdinv5
+ dout_5 dout_6 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_5_0
+ dout_6 n_5_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_5_1
+ dout_6 n_5_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_5_2
+ dout_6 n_5_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_5_3
+ dout_6 n_5_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdinv6
+ dout_6 dout_7 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_6_0
+ dout_7 n_6_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_6_1
+ dout_7 n_6_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_6_2
+ dout_7 n_6_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_6_3
+ dout_7 n_6_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdinv7
+ dout_7 dout_8 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_7_0
+ dout_8 n_7_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_7_1
+ dout_8 n_7_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_7_2
+ dout_8 n_7_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_7_3
+ dout_8 n_7_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdinv8
+ dout_8 out vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_8_0
+ out n_8_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_8_1
+ out n_8_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_8_2
+ out n_8_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
Xdload_8_3
+ out n_8_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_20
.ENDS sky130_sram_1kbyte_1rw_32x256_8_delay_chain

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pnand3
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpnand3_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand3_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand3_pmos3 Z C vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand3_nmos1 Z C net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand3_nmos2 net1 B net2 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand3_nmos3 net2 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pnand3

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=9 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=9 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_14
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 40
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=9 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=9 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_14

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pdriver_4
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [40]
Xbuf_inv1
+ A Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_14
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pdriver_4

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pand3
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 40
Xpand3_nand
+ A B C zb_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pnand3
Xpand3_inv
+ zb_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pdriver_4
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pand3

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_16
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_16

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=8 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=8 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_15
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 33
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=8 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=8 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_15

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pdriver_5
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [33]
Xbuf_inv1
+ A Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_15
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pdriver_5

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pand3_0
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 33
Xpand3_nand
+ A B C zb_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pnand3
Xpand3_inv
+ zb_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pdriver_5
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pand3_0

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pnand2
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpnand2_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_nmos1 Z B net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand2_nmos2 net1 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pnand2

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=3 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=3 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_4
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 12
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=3 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=3 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_4

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pdriver_1
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [12]
Xbuf_inv1
+ A Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_4
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pdriver_1

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pand2_1
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 12
Xpand2_nand
+ A B zb_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pnand2
Xpand2_inv
+ zb_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pdriver_1
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pand2_1

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=10 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=10 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_19
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 43
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=10 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=10 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_19

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=6 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=6 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_18
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 14
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=6 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=6 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_18

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=2 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 2.0
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=2 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=2 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_17
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 5
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=2 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=2 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_17

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pdriver_6
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 2, 5, 14, 43]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_7
Xbuf_inv2
+ Zb1_int Zb2_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_7
Xbuf_inv3
+ Zb2_int Zb3_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv
Xbuf_inv4
+ Zb3_int Zb4_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_17
Xbuf_inv5
+ Zb4_int Zb5_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_18
Xbuf_inv6
+ Zb5_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_19
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pdriver_6

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=5 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=5 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_13
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 21
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=5 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=5 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_13

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_12
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 7
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_12

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pdriver_3
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [7, 21]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_12
Xbuf_inv2
+ Zb1_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_13
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pdriver_3

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_3
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 4
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_3
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* SPICE3 file created from sky130_fd_bd_sram__openram_dff.ext - technology: EFS8A

.subckt sky130_fd_bd_sram__openram_dff D Q CLK VDD GND
X1000 a_511_725# a_n8_115# VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1001 a_353_115# CLK a_11_624# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1002 a_353_725# a_203_89# a_11_624# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1003 a_11_624# a_203_89# a_161_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1004 a_11_624# CLK a_161_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1005 GND Q a_703_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1006 VDD Q a_703_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1007 a_203_89# CLK GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1008 a_203_89# CLK VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1009 a_161_115# D GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1010 a_161_725# D VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1011 GND a_11_624# a_n8_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1012 a_703_115# a_203_89# ON GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1013 VDD a_11_624# a_n8_115# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1014 a_703_725# CLK ON VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1015 Q ON VDD VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1016 Q ON GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1017 ON a_203_89# a_511_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1018 ON CLK a_511_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1019 GND a_n8_115# a_353_115# GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X1020 VDD a_n8_115# a_353_725# VDD sky130_fd_pr__pfet_01v8 W=3 L=0.15
X1021 a_511_115# a_n8_115# GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
.ends

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_2
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 2
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=2 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_2

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_dff_buf_0
+ D Q Qb clk vdd gnd
* INPUT : D 
* OUTPUT: Q 
* OUTPUT: Qb 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_buf_dff
+ D qint clk vdd gnd
+ sky130_fd_bd_sram__openram_dff
Xdff_buf_inv1
+ qint Qb vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_2
Xdff_buf_inv2
+ Qb Q vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_3
.ENDS sky130_sram_1kbyte_1rw_32x256_8_dff_buf_0

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_dff_buf_array
+ din_0 din_1 dout_0 dout_bar_0 dout_1 dout_bar_1 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_bar_0 
* OUTPUT: dout_1 
* OUTPUT: dout_bar_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 2 cols: 1
* inv1: 2 inv2: 4
Xdff_r0_c0
+ din_0 dout_0 dout_bar_0 clk vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_dff_buf_0
Xdff_r1_c0
+ din_1 dout_1 dout_bar_1 clk vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_dff_buf_0
.ENDS sky130_sram_1kbyte_1rw_32x256_8_dff_buf_array

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_control_logic_rw
+ csb web clk rbl_bl s_en w_en p_en_bar wl_en clk_buf vdd gnd
* INPUT : csb 
* INPUT : web 
* INPUT : clk 
* INPUT : rbl_bl 
* OUTPUT: s_en 
* OUTPUT: w_en 
* OUTPUT: p_en_bar 
* OUTPUT: wl_en 
* OUTPUT: clk_buf 
* POWER : vdd 
* GROUND: gnd 
* num_rows: 65
* words_per_row: 4
* word_size 32
Xctrl_dffs
+ csb web cs_bar cs we_bar we clk_buf vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_dff_buf_array
Xclkbuf
+ clk clk_buf vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pdriver_2
Xinv_clk_bar
+ clk_buf clk_bar vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_16
Xand2_gated_clk_bar
+ clk_bar cs gated_clk_bar vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand2_1
Xand2_gated_clk_buf
+ clk_buf cs gated_clk_buf vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand2_1
Xbuf_wl_en
+ gated_clk_bar wl_en vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pdriver_3
Xrbl_bl_delay_inv
+ rbl_bl_delay rbl_bl_delay_bar vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_16
Xw_en_and
+ we rbl_bl_delay_bar gated_clk_bar w_en vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand3
Xbuf_s_en_and
+ rbl_bl_delay gated_clk_bar we_bar s_en vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand3_0
Xdelay_chain
+ rbl_bl rbl_bl_delay vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_delay_chain
Xnand_p_en_bar
+ gated_clk_buf rbl_bl_delay p_en_bar_unbuf vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pnand2_1
Xbuf_p_en_bar
+ p_en_bar_unbuf p_en_bar vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pdriver_6
.ENDS sky130_sram_1kbyte_1rw_32x256_8_control_logic_rw

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_wmask_dff
+ din_0 din_1 din_2 din_3 dout_0 dout_1 dout_2 dout_3 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 4
Xdff_r0_c0
+ din_0 dout_0 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c1
+ din_1 dout_1 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c2
+ din_2 dout_2 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c3
+ din_3 dout_3 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
.ENDS sky130_sram_1kbyte_1rw_32x256_8_wmask_dff

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_spare_wen_dff
+ din_0 dout_0 clk vdd gnd
* INPUT : din_0 
* OUTPUT: dout_0 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 1
Xdff_r0_c0
+ din_0 dout_0 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
.ENDS sky130_sram_1kbyte_1rw_32x256_8_spare_wen_dff

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_col_addr_dff
+ din_0 din_1 dout_0 dout_1 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 2
Xdff_r0_c0
+ din_0 dout_0 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c1
+ din_1 dout_1 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
.ENDS sky130_sram_1kbyte_1rw_32x256_8_col_addr_dff

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_1
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_1

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_0

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pdriver_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1]
Xbuf_inv1
+ A Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_0
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pdriver_0

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pnand2_0
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpnand2_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_nmos1 Z B net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand2_nmos2 net1 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pnand2_0

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pand2_0
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand2_nand
+ A B zb_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pnand2_0
Xpand2_inv
+ zb_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pdriver_0
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pand2_0

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_hierarchical_predecode2x4_0
+ in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0
+ in_0 inbar_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_1
Xpre_inv_1
+ in_1 inbar_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_1
XXpre2x4_and_0
+ inbar_0 inbar_1 out_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand2_0
XXpre2x4_and_1
+ in_0 inbar_1 out_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand2_0
XXpre2x4_and_2
+ inbar_0 in_1 out_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand2_0
XXpre2x4_and_3
+ in_0 in_1 out_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand2_0
.ENDS sky130_sram_1kbyte_1rw_32x256_8_hierarchical_predecode2x4_0

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_column_decoder
+ in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xcolumn_decoder
+ in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_hierarchical_predecode2x4_0
.ENDS sky130_sram_1kbyte_1rw_32x256_8_column_decoder
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

*********************** "sky130_fd_bd_sram__openram_sense_amp" ******************************

.SUBCKT sky130_fd_bd_sram__openram_sense_amp BL BR DOUT EN VDD GND
X1000 GND EN a_56_432# GND sky130_fd_pr__nfet_01v8 W=0.65 L=0.15
X1001 a_56_432# dint_bar dint GND sky130_fd_pr__nfet_01v8 W=0.65 L=0.15
X1002 dint_bar dint a_56_432# GND sky130_fd_pr__nfet_01v8 W=0.65 L=0.15

X1003 VDD dint_bar dint VDD sky130_fd_pr__pfet_01v8 W=1.26 L=0.15
X1004 dint_bar dint VDD VDD sky130_fd_pr__pfet_01v8 W=1.26 L=0.15

X1005 BL EN dint VDD sky130_fd_pr__pfet_01v8 W=2 L=0.15
X1006 dint_bar EN BR VDD sky130_fd_pr__pfet_01v8 W=2 L=0.15

X1007 VDD dint_bar DOUT VDD sky130_fd_pr__pfet_01v8 W=1.26 L=0.15
X1008 DOUT dint_bar GND GND sky130_fd_pr__nfet_01v8 W=0.65 L=0.15

.ENDS sky130_fd_bd_sram__openram_sense_amp

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_sense_amp_array
+ data_0 bl_0 br_0 data_1 bl_1 br_1 data_2 bl_2 br_2 data_3 bl_3 br_3
+ data_4 bl_4 br_4 data_5 bl_5 br_5 data_6 bl_6 br_6 data_7 bl_7 br_7
+ data_8 bl_8 br_8 data_9 bl_9 br_9 data_10 bl_10 br_10 data_11 bl_11
+ br_11 data_12 bl_12 br_12 data_13 bl_13 br_13 data_14 bl_14 br_14
+ data_15 bl_15 br_15 data_16 bl_16 br_16 data_17 bl_17 br_17 data_18
+ bl_18 br_18 data_19 bl_19 br_19 data_20 bl_20 br_20 data_21 bl_21
+ br_21 data_22 bl_22 br_22 data_23 bl_23 br_23 data_24 bl_24 br_24
+ data_25 bl_25 br_25 data_26 bl_26 br_26 data_27 bl_27 br_27 data_28
+ bl_28 br_28 data_29 bl_29 br_29 data_30 bl_30 br_30 data_31 bl_31
+ br_31 data_32 bl_32 br_32 en vdd gnd
* OUTPUT: data_0 
* INPUT : bl_0 
* INPUT : br_0 
* OUTPUT: data_1 
* INPUT : bl_1 
* INPUT : br_1 
* OUTPUT: data_2 
* INPUT : bl_2 
* INPUT : br_2 
* OUTPUT: data_3 
* INPUT : bl_3 
* INPUT : br_3 
* OUTPUT: data_4 
* INPUT : bl_4 
* INPUT : br_4 
* OUTPUT: data_5 
* INPUT : bl_5 
* INPUT : br_5 
* OUTPUT: data_6 
* INPUT : bl_6 
* INPUT : br_6 
* OUTPUT: data_7 
* INPUT : bl_7 
* INPUT : br_7 
* OUTPUT: data_8 
* INPUT : bl_8 
* INPUT : br_8 
* OUTPUT: data_9 
* INPUT : bl_9 
* INPUT : br_9 
* OUTPUT: data_10 
* INPUT : bl_10 
* INPUT : br_10 
* OUTPUT: data_11 
* INPUT : bl_11 
* INPUT : br_11 
* OUTPUT: data_12 
* INPUT : bl_12 
* INPUT : br_12 
* OUTPUT: data_13 
* INPUT : bl_13 
* INPUT : br_13 
* OUTPUT: data_14 
* INPUT : bl_14 
* INPUT : br_14 
* OUTPUT: data_15 
* INPUT : bl_15 
* INPUT : br_15 
* OUTPUT: data_16 
* INPUT : bl_16 
* INPUT : br_16 
* OUTPUT: data_17 
* INPUT : bl_17 
* INPUT : br_17 
* OUTPUT: data_18 
* INPUT : bl_18 
* INPUT : br_18 
* OUTPUT: data_19 
* INPUT : bl_19 
* INPUT : br_19 
* OUTPUT: data_20 
* INPUT : bl_20 
* INPUT : br_20 
* OUTPUT: data_21 
* INPUT : bl_21 
* INPUT : br_21 
* OUTPUT: data_22 
* INPUT : bl_22 
* INPUT : br_22 
* OUTPUT: data_23 
* INPUT : bl_23 
* INPUT : br_23 
* OUTPUT: data_24 
* INPUT : bl_24 
* INPUT : br_24 
* OUTPUT: data_25 
* INPUT : bl_25 
* INPUT : br_25 
* OUTPUT: data_26 
* INPUT : bl_26 
* INPUT : br_26 
* OUTPUT: data_27 
* INPUT : bl_27 
* INPUT : br_27 
* OUTPUT: data_28 
* INPUT : bl_28 
* INPUT : br_28 
* OUTPUT: data_29 
* INPUT : bl_29 
* INPUT : br_29 
* OUTPUT: data_30 
* INPUT : bl_30 
* INPUT : br_30 
* OUTPUT: data_31 
* INPUT : bl_31 
* INPUT : br_31 
* OUTPUT: data_32 
* INPUT : bl_32 
* INPUT : br_32 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* word_size 32
* words_per_row: 4
Xsa_d0
+ bl_0 br_0 data_0 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d1
+ bl_1 br_1 data_1 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d2
+ bl_2 br_2 data_2 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d3
+ bl_3 br_3 data_3 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d4
+ bl_4 br_4 data_4 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d5
+ bl_5 br_5 data_5 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d6
+ bl_6 br_6 data_6 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d7
+ bl_7 br_7 data_7 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d8
+ bl_8 br_8 data_8 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d9
+ bl_9 br_9 data_9 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d10
+ bl_10 br_10 data_10 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d11
+ bl_11 br_11 data_11 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d12
+ bl_12 br_12 data_12 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d13
+ bl_13 br_13 data_13 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d14
+ bl_14 br_14 data_14 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d15
+ bl_15 br_15 data_15 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d16
+ bl_16 br_16 data_16 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d17
+ bl_17 br_17 data_17 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d18
+ bl_18 br_18 data_18 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d19
+ bl_19 br_19 data_19 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d20
+ bl_20 br_20 data_20 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d21
+ bl_21 br_21 data_21 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d22
+ bl_22 br_22 data_22 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d23
+ bl_23 br_23 data_23 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d24
+ bl_24 br_24 data_24 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d25
+ bl_25 br_25 data_25 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d26
+ bl_26 br_26 data_26 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d27
+ bl_27 br_27 data_27 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d28
+ bl_28 br_28 data_28 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d29
+ bl_29 br_29 data_29 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d30
+ bl_30 br_30 data_30 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d31
+ bl_31 br_31 data_31 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
Xsa_d32
+ bl_32 br_32 data_32 en vdd gnd
+ sky130_fd_bd_sram__openram_sense_amp
.ENDS sky130_sram_1kbyte_1rw_32x256_8_sense_amp_array
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

*********************** "sky130_fd_bd_sram__openram_write_driver" ******************************

.SUBCKT sky130_fd_bd_sram__openram_write_driver DIN BL BR EN VDD GND

**** Inverter to conver Data_in to data_in_bar ******
* din_bar = inv(DIN)
X_1 din_bar DIN GND GND sky130_fd_pr__nfet_01v8 W=0.36 L=0.15
X_2 din_bar DIN VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15

**** 2input nand gate follwed by inverter to drive BL ******
* din_bar_gated = nand(EN, DIN)
X_3 din_bar_gated EN net_7 GND sky130_fd_pr__nfet_01v8 W=0.55 L=0.15
X_4 net_7 DIN GND GND sky130_fd_pr__nfet_01v8 W=0.55 L=0.15
X_5 din_bar_gated EN VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
X_6 din_bar_gated DIN VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
* din_bar_gated_bar = inv(din_bar_gated)
X_7 din_bar_gated_bar din_bar_gated VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
X_8 din_bar_gated_bar din_bar_gated GND GND sky130_fd_pr__nfet_01v8 W=0.36 L=0.15

**** 2input nand gate follwed by inverter to drive BR******
* din_gated = nand(EN, din_bar)
X_9 din_gated EN VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
X_10 din_gated EN net_8 GND sky130_fd_pr__nfet_01v8 W=0.55 L=0.15
X_11 net_8 din_bar GND GND sky130_fd_pr__nfet_01v8 W=0.55 L=0.15
X_12 din_gated din_bar VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
* din_gated_bar = inv(din_gated)
X_13 din_gated_bar din_gated VDD VDD sky130_fd_pr__pfet_01v8 W=0.55 L=0.15
X_14 din_gated_bar din_gated GND GND sky130_fd_pr__nfet_01v8 W=0.36 L=0.15

************************************************
* pull down with EN enable
X_15 BL din_gated_bar GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15
X_16 BR din_bar_gated_bar GND GND sky130_fd_pr__nfet_01v8 W=1 L=0.15

.ENDS sky130_fd_bd_sram__openram_write_driver

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_write_driver_array
+ data_0 data_1 data_2 data_3 data_4 data_5 data_6 data_7 data_8 data_9
+ data_10 data_11 data_12 data_13 data_14 data_15 data_16 data_17
+ data_18 data_19 data_20 data_21 data_22 data_23 data_24 data_25
+ data_26 data_27 data_28 data_29 data_30 data_31 data_32 bl_0 br_0 bl_1
+ br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8
+ br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14
+ br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19
+ bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25
+ br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30
+ bl_31 br_31 bl_32 br_32 en_0 en_1 en_2 en_3 en_4 vdd gnd
* INPUT : data_0 
* INPUT : data_1 
* INPUT : data_2 
* INPUT : data_3 
* INPUT : data_4 
* INPUT : data_5 
* INPUT : data_6 
* INPUT : data_7 
* INPUT : data_8 
* INPUT : data_9 
* INPUT : data_10 
* INPUT : data_11 
* INPUT : data_12 
* INPUT : data_13 
* INPUT : data_14 
* INPUT : data_15 
* INPUT : data_16 
* INPUT : data_17 
* INPUT : data_18 
* INPUT : data_19 
* INPUT : data_20 
* INPUT : data_21 
* INPUT : data_22 
* INPUT : data_23 
* INPUT : data_24 
* INPUT : data_25 
* INPUT : data_26 
* INPUT : data_27 
* INPUT : data_28 
* INPUT : data_29 
* INPUT : data_30 
* INPUT : data_31 
* INPUT : data_32 
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* INPUT : en_0 
* INPUT : en_1 
* INPUT : en_2 
* INPUT : en_3 
* INPUT : en_4 
* POWER : vdd 
* GROUND: gnd 
* columns: 128
* word_size 32
Xwrite_driver0
+ data_0 bl_0 br_0 en_0 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver4
+ data_1 bl_1 br_1 en_0 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver8
+ data_2 bl_2 br_2 en_0 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver12
+ data_3 bl_3 br_3 en_0 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver16
+ data_4 bl_4 br_4 en_0 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver20
+ data_5 bl_5 br_5 en_0 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver24
+ data_6 bl_6 br_6 en_0 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver28
+ data_7 bl_7 br_7 en_0 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver32
+ data_8 bl_8 br_8 en_1 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver36
+ data_9 bl_9 br_9 en_1 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver40
+ data_10 bl_10 br_10 en_1 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver44
+ data_11 bl_11 br_11 en_1 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver48
+ data_12 bl_12 br_12 en_1 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver52
+ data_13 bl_13 br_13 en_1 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver56
+ data_14 bl_14 br_14 en_1 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver60
+ data_15 bl_15 br_15 en_1 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver64
+ data_16 bl_16 br_16 en_2 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver68
+ data_17 bl_17 br_17 en_2 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver72
+ data_18 bl_18 br_18 en_2 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver76
+ data_19 bl_19 br_19 en_2 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver80
+ data_20 bl_20 br_20 en_2 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver84
+ data_21 bl_21 br_21 en_2 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver88
+ data_22 bl_22 br_22 en_2 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver92
+ data_23 bl_23 br_23 en_2 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver96
+ data_24 bl_24 br_24 en_3 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver100
+ data_25 bl_25 br_25 en_3 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver104
+ data_26 bl_26 br_26 en_3 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver108
+ data_27 bl_27 br_27 en_3 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver112
+ data_28 bl_28 br_28 en_3 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver116
+ data_29 bl_29 br_29 en_3 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver120
+ data_30 bl_30 br_30 en_3 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver124
+ data_31 bl_31 br_31 en_3 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
Xwrite_driver128
+ data_32 bl_32 br_32 en_4 vdd gnd
+ sky130_fd_bd_sram__openram_write_driver
.ENDS sky130_sram_1kbyte_1rw_32x256_8_write_driver_array

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pdriver
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [2.0]
Xbuf_inv1
+ A Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pdriver

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pand2
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 2.0
Xpand2_nand
+ A B zb_int vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pnand2
Xpand2_inv
+ zb_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pdriver
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pand2

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_write_mask_and_array
+ wmask_in_0 wmask_in_1 wmask_in_2 wmask_in_3 en wmask_out_0 wmask_out_1
+ wmask_out_2 wmask_out_3 vdd gnd
* INPUT : wmask_in_0 
* INPUT : wmask_in_1 
* INPUT : wmask_in_2 
* INPUT : wmask_in_3 
* INPUT : en 
* OUTPUT: wmask_out_0 
* OUTPUT: wmask_out_1 
* OUTPUT: wmask_out_2 
* OUTPUT: wmask_out_3 
* POWER : vdd 
* GROUND: gnd 
* columns: 128
* word_size 32
* write_size 8
Xand2_0
+ wmask_in_0 en wmask_out_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand2
Xand2_1
+ wmask_in_1 en wmask_out_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand2
Xand2_2
+ wmask_in_2 en wmask_out_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand2
Xand2_3
+ wmask_in_3 en wmask_out_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pand2
.ENDS sky130_sram_1kbyte_1rw_32x256_8_write_mask_and_array

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.88 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_column_mux
+ bl br bl_out br_out sel gnd
* INOUT : bl 
* INOUT : br 
* INOUT : bl_out 
* INOUT : br_out 
* INOUT : sel 
* INOUT : gnd 
Xmux_tx1 bl sel bl_out gnd sky130_fd_pr__nfet_01v8 m=1 w=2.88 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u
Xmux_tx2 br sel br_out gnd sky130_fd_pr__nfet_01v8 m=1 w=2.88 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_column_mux

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_column_mux_array
+ bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18
+ br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23
+ bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34
+ bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40
+ br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51
+ br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67
+ bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73
+ br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78
+ bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84
+ br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89
+ bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95
+ br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100
+ bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105
+ bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110
+ bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115
+ bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120
+ bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125
+ bl_126 br_126 bl_127 br_127 sel_0 sel_1 sel_2 sel_3 bl_out_0 br_out_0
+ bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4
+ br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7
+ bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11
+ br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14
+ bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18
+ br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21
+ bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25
+ br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28
+ bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : sel_0 
* INOUT : sel_1 
* INOUT : sel_2 
* INOUT : sel_3 
* INOUT : bl_out_0 
* INOUT : br_out_0 
* INOUT : bl_out_1 
* INOUT : br_out_1 
* INOUT : bl_out_2 
* INOUT : br_out_2 
* INOUT : bl_out_3 
* INOUT : br_out_3 
* INOUT : bl_out_4 
* INOUT : br_out_4 
* INOUT : bl_out_5 
* INOUT : br_out_5 
* INOUT : bl_out_6 
* INOUT : br_out_6 
* INOUT : bl_out_7 
* INOUT : br_out_7 
* INOUT : bl_out_8 
* INOUT : br_out_8 
* INOUT : bl_out_9 
* INOUT : br_out_9 
* INOUT : bl_out_10 
* INOUT : br_out_10 
* INOUT : bl_out_11 
* INOUT : br_out_11 
* INOUT : bl_out_12 
* INOUT : br_out_12 
* INOUT : bl_out_13 
* INOUT : br_out_13 
* INOUT : bl_out_14 
* INOUT : br_out_14 
* INOUT : bl_out_15 
* INOUT : br_out_15 
* INOUT : bl_out_16 
* INOUT : br_out_16 
* INOUT : bl_out_17 
* INOUT : br_out_17 
* INOUT : bl_out_18 
* INOUT : br_out_18 
* INOUT : bl_out_19 
* INOUT : br_out_19 
* INOUT : bl_out_20 
* INOUT : br_out_20 
* INOUT : bl_out_21 
* INOUT : br_out_21 
* INOUT : bl_out_22 
* INOUT : br_out_22 
* INOUT : bl_out_23 
* INOUT : br_out_23 
* INOUT : bl_out_24 
* INOUT : br_out_24 
* INOUT : bl_out_25 
* INOUT : br_out_25 
* INOUT : bl_out_26 
* INOUT : br_out_26 
* INOUT : bl_out_27 
* INOUT : br_out_27 
* INOUT : bl_out_28 
* INOUT : br_out_28 
* INOUT : bl_out_29 
* INOUT : br_out_29 
* INOUT : bl_out_30 
* INOUT : br_out_30 
* INOUT : bl_out_31 
* INOUT : br_out_31 
* INOUT : gnd 
* cols: 128 word_size: 32 bl: bl br: br
XXMUX0
+ bl_0 br_0 bl_out_0 br_out_0 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX1
+ bl_1 br_1 bl_out_0 br_out_0 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX2
+ bl_2 br_2 bl_out_0 br_out_0 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX3
+ bl_3 br_3 bl_out_0 br_out_0 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX4
+ bl_4 br_4 bl_out_1 br_out_1 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX5
+ bl_5 br_5 bl_out_1 br_out_1 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX6
+ bl_6 br_6 bl_out_1 br_out_1 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX7
+ bl_7 br_7 bl_out_1 br_out_1 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX8
+ bl_8 br_8 bl_out_2 br_out_2 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX9
+ bl_9 br_9 bl_out_2 br_out_2 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX10
+ bl_10 br_10 bl_out_2 br_out_2 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX11
+ bl_11 br_11 bl_out_2 br_out_2 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX12
+ bl_12 br_12 bl_out_3 br_out_3 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX13
+ bl_13 br_13 bl_out_3 br_out_3 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX14
+ bl_14 br_14 bl_out_3 br_out_3 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX15
+ bl_15 br_15 bl_out_3 br_out_3 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX16
+ bl_16 br_16 bl_out_4 br_out_4 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX17
+ bl_17 br_17 bl_out_4 br_out_4 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX18
+ bl_18 br_18 bl_out_4 br_out_4 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX19
+ bl_19 br_19 bl_out_4 br_out_4 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX20
+ bl_20 br_20 bl_out_5 br_out_5 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX21
+ bl_21 br_21 bl_out_5 br_out_5 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX22
+ bl_22 br_22 bl_out_5 br_out_5 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX23
+ bl_23 br_23 bl_out_5 br_out_5 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX24
+ bl_24 br_24 bl_out_6 br_out_6 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX25
+ bl_25 br_25 bl_out_6 br_out_6 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX26
+ bl_26 br_26 bl_out_6 br_out_6 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX27
+ bl_27 br_27 bl_out_6 br_out_6 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX28
+ bl_28 br_28 bl_out_7 br_out_7 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX29
+ bl_29 br_29 bl_out_7 br_out_7 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX30
+ bl_30 br_30 bl_out_7 br_out_7 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX31
+ bl_31 br_31 bl_out_7 br_out_7 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX32
+ bl_32 br_32 bl_out_8 br_out_8 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX33
+ bl_33 br_33 bl_out_8 br_out_8 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX34
+ bl_34 br_34 bl_out_8 br_out_8 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX35
+ bl_35 br_35 bl_out_8 br_out_8 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX36
+ bl_36 br_36 bl_out_9 br_out_9 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX37
+ bl_37 br_37 bl_out_9 br_out_9 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX38
+ bl_38 br_38 bl_out_9 br_out_9 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX39
+ bl_39 br_39 bl_out_9 br_out_9 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX40
+ bl_40 br_40 bl_out_10 br_out_10 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX41
+ bl_41 br_41 bl_out_10 br_out_10 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX42
+ bl_42 br_42 bl_out_10 br_out_10 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX43
+ bl_43 br_43 bl_out_10 br_out_10 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX44
+ bl_44 br_44 bl_out_11 br_out_11 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX45
+ bl_45 br_45 bl_out_11 br_out_11 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX46
+ bl_46 br_46 bl_out_11 br_out_11 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX47
+ bl_47 br_47 bl_out_11 br_out_11 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX48
+ bl_48 br_48 bl_out_12 br_out_12 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX49
+ bl_49 br_49 bl_out_12 br_out_12 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX50
+ bl_50 br_50 bl_out_12 br_out_12 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX51
+ bl_51 br_51 bl_out_12 br_out_12 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX52
+ bl_52 br_52 bl_out_13 br_out_13 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX53
+ bl_53 br_53 bl_out_13 br_out_13 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX54
+ bl_54 br_54 bl_out_13 br_out_13 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX55
+ bl_55 br_55 bl_out_13 br_out_13 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX56
+ bl_56 br_56 bl_out_14 br_out_14 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX57
+ bl_57 br_57 bl_out_14 br_out_14 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX58
+ bl_58 br_58 bl_out_14 br_out_14 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX59
+ bl_59 br_59 bl_out_14 br_out_14 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX60
+ bl_60 br_60 bl_out_15 br_out_15 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX61
+ bl_61 br_61 bl_out_15 br_out_15 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX62
+ bl_62 br_62 bl_out_15 br_out_15 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX63
+ bl_63 br_63 bl_out_15 br_out_15 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX64
+ bl_64 br_64 bl_out_16 br_out_16 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX65
+ bl_65 br_65 bl_out_16 br_out_16 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX66
+ bl_66 br_66 bl_out_16 br_out_16 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX67
+ bl_67 br_67 bl_out_16 br_out_16 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX68
+ bl_68 br_68 bl_out_17 br_out_17 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX69
+ bl_69 br_69 bl_out_17 br_out_17 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX70
+ bl_70 br_70 bl_out_17 br_out_17 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX71
+ bl_71 br_71 bl_out_17 br_out_17 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX72
+ bl_72 br_72 bl_out_18 br_out_18 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX73
+ bl_73 br_73 bl_out_18 br_out_18 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX74
+ bl_74 br_74 bl_out_18 br_out_18 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX75
+ bl_75 br_75 bl_out_18 br_out_18 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX76
+ bl_76 br_76 bl_out_19 br_out_19 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX77
+ bl_77 br_77 bl_out_19 br_out_19 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX78
+ bl_78 br_78 bl_out_19 br_out_19 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX79
+ bl_79 br_79 bl_out_19 br_out_19 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX80
+ bl_80 br_80 bl_out_20 br_out_20 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX81
+ bl_81 br_81 bl_out_20 br_out_20 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX82
+ bl_82 br_82 bl_out_20 br_out_20 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX83
+ bl_83 br_83 bl_out_20 br_out_20 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX84
+ bl_84 br_84 bl_out_21 br_out_21 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX85
+ bl_85 br_85 bl_out_21 br_out_21 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX86
+ bl_86 br_86 bl_out_21 br_out_21 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX87
+ bl_87 br_87 bl_out_21 br_out_21 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX88
+ bl_88 br_88 bl_out_22 br_out_22 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX89
+ bl_89 br_89 bl_out_22 br_out_22 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX90
+ bl_90 br_90 bl_out_22 br_out_22 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX91
+ bl_91 br_91 bl_out_22 br_out_22 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX92
+ bl_92 br_92 bl_out_23 br_out_23 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX93
+ bl_93 br_93 bl_out_23 br_out_23 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX94
+ bl_94 br_94 bl_out_23 br_out_23 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX95
+ bl_95 br_95 bl_out_23 br_out_23 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX96
+ bl_96 br_96 bl_out_24 br_out_24 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX97
+ bl_97 br_97 bl_out_24 br_out_24 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX98
+ bl_98 br_98 bl_out_24 br_out_24 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX99
+ bl_99 br_99 bl_out_24 br_out_24 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX100
+ bl_100 br_100 bl_out_25 br_out_25 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX101
+ bl_101 br_101 bl_out_25 br_out_25 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX102
+ bl_102 br_102 bl_out_25 br_out_25 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX103
+ bl_103 br_103 bl_out_25 br_out_25 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX104
+ bl_104 br_104 bl_out_26 br_out_26 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX105
+ bl_105 br_105 bl_out_26 br_out_26 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX106
+ bl_106 br_106 bl_out_26 br_out_26 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX107
+ bl_107 br_107 bl_out_26 br_out_26 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX108
+ bl_108 br_108 bl_out_27 br_out_27 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX109
+ bl_109 br_109 bl_out_27 br_out_27 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX110
+ bl_110 br_110 bl_out_27 br_out_27 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX111
+ bl_111 br_111 bl_out_27 br_out_27 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX112
+ bl_112 br_112 bl_out_28 br_out_28 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX113
+ bl_113 br_113 bl_out_28 br_out_28 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX114
+ bl_114 br_114 bl_out_28 br_out_28 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX115
+ bl_115 br_115 bl_out_28 br_out_28 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX116
+ bl_116 br_116 bl_out_29 br_out_29 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX117
+ bl_117 br_117 bl_out_29 br_out_29 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX118
+ bl_118 br_118 bl_out_29 br_out_29 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX119
+ bl_119 br_119 bl_out_29 br_out_29 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX120
+ bl_120 br_120 bl_out_30 br_out_30 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX121
+ bl_121 br_121 bl_out_30 br_out_30 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX122
+ bl_122 br_122 bl_out_30 br_out_30 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX123
+ bl_123 br_123 bl_out_30 br_out_30 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX124
+ bl_124 br_124 bl_out_31 br_out_31 sel_0 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX125
+ bl_125 br_125 bl_out_31 br_out_31 sel_1 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX126
+ bl_126 br_126 bl_out_31 br_out_31 sel_2 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
XXMUX127
+ bl_127 br_127 bl_out_31 br_out_31 sel_3 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux
.ENDS sky130_sram_1kbyte_1rw_32x256_8_column_mux_array

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_precharge_0
+ bl br en_bar vdd
* OUTPUT: bl 
* OUTPUT: br 
* INPUT : en_bar 
* POWER : vdd 
Xlower_pmos bl en_bar br vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
Xupper_pmos1 bl en_bar vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
Xupper_pmos2 br en_bar vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=0.15 pd=1.40 ps=1.40 as=0.21u ad=0.21u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_precharge_0

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_precharge_array
+ bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18
+ br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23
+ bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34
+ bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40
+ br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51
+ br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67
+ bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73
+ br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78
+ bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84
+ br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89
+ bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95
+ br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100
+ bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105
+ bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110
+ bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115
+ bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120
+ bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125
+ bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 en_bar vdd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* OUTPUT: bl_65 
* OUTPUT: br_65 
* OUTPUT: bl_66 
* OUTPUT: br_66 
* OUTPUT: bl_67 
* OUTPUT: br_67 
* OUTPUT: bl_68 
* OUTPUT: br_68 
* OUTPUT: bl_69 
* OUTPUT: br_69 
* OUTPUT: bl_70 
* OUTPUT: br_70 
* OUTPUT: bl_71 
* OUTPUT: br_71 
* OUTPUT: bl_72 
* OUTPUT: br_72 
* OUTPUT: bl_73 
* OUTPUT: br_73 
* OUTPUT: bl_74 
* OUTPUT: br_74 
* OUTPUT: bl_75 
* OUTPUT: br_75 
* OUTPUT: bl_76 
* OUTPUT: br_76 
* OUTPUT: bl_77 
* OUTPUT: br_77 
* OUTPUT: bl_78 
* OUTPUT: br_78 
* OUTPUT: bl_79 
* OUTPUT: br_79 
* OUTPUT: bl_80 
* OUTPUT: br_80 
* OUTPUT: bl_81 
* OUTPUT: br_81 
* OUTPUT: bl_82 
* OUTPUT: br_82 
* OUTPUT: bl_83 
* OUTPUT: br_83 
* OUTPUT: bl_84 
* OUTPUT: br_84 
* OUTPUT: bl_85 
* OUTPUT: br_85 
* OUTPUT: bl_86 
* OUTPUT: br_86 
* OUTPUT: bl_87 
* OUTPUT: br_87 
* OUTPUT: bl_88 
* OUTPUT: br_88 
* OUTPUT: bl_89 
* OUTPUT: br_89 
* OUTPUT: bl_90 
* OUTPUT: br_90 
* OUTPUT: bl_91 
* OUTPUT: br_91 
* OUTPUT: bl_92 
* OUTPUT: br_92 
* OUTPUT: bl_93 
* OUTPUT: br_93 
* OUTPUT: bl_94 
* OUTPUT: br_94 
* OUTPUT: bl_95 
* OUTPUT: br_95 
* OUTPUT: bl_96 
* OUTPUT: br_96 
* OUTPUT: bl_97 
* OUTPUT: br_97 
* OUTPUT: bl_98 
* OUTPUT: br_98 
* OUTPUT: bl_99 
* OUTPUT: br_99 
* OUTPUT: bl_100 
* OUTPUT: br_100 
* OUTPUT: bl_101 
* OUTPUT: br_101 
* OUTPUT: bl_102 
* OUTPUT: br_102 
* OUTPUT: bl_103 
* OUTPUT: br_103 
* OUTPUT: bl_104 
* OUTPUT: br_104 
* OUTPUT: bl_105 
* OUTPUT: br_105 
* OUTPUT: bl_106 
* OUTPUT: br_106 
* OUTPUT: bl_107 
* OUTPUT: br_107 
* OUTPUT: bl_108 
* OUTPUT: br_108 
* OUTPUT: bl_109 
* OUTPUT: br_109 
* OUTPUT: bl_110 
* OUTPUT: br_110 
* OUTPUT: bl_111 
* OUTPUT: br_111 
* OUTPUT: bl_112 
* OUTPUT: br_112 
* OUTPUT: bl_113 
* OUTPUT: br_113 
* OUTPUT: bl_114 
* OUTPUT: br_114 
* OUTPUT: bl_115 
* OUTPUT: br_115 
* OUTPUT: bl_116 
* OUTPUT: br_116 
* OUTPUT: bl_117 
* OUTPUT: br_117 
* OUTPUT: bl_118 
* OUTPUT: br_118 
* OUTPUT: bl_119 
* OUTPUT: br_119 
* OUTPUT: bl_120 
* OUTPUT: br_120 
* OUTPUT: bl_121 
* OUTPUT: br_121 
* OUTPUT: bl_122 
* OUTPUT: br_122 
* OUTPUT: bl_123 
* OUTPUT: br_123 
* OUTPUT: bl_124 
* OUTPUT: br_124 
* OUTPUT: bl_125 
* OUTPUT: br_125 
* OUTPUT: bl_126 
* OUTPUT: br_126 
* OUTPUT: bl_127 
* OUTPUT: br_127 
* OUTPUT: bl_128 
* OUTPUT: br_128 
* OUTPUT: bl_129 
* OUTPUT: br_129 
* INPUT : en_bar 
* POWER : vdd 
* cols: 130 size: 1 bl: bl br: br
Xpre_column_0
+ bl_0 br_0 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_1
+ bl_1 br_1 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_2
+ bl_2 br_2 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_3
+ bl_3 br_3 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_4
+ bl_4 br_4 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_5
+ bl_5 br_5 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_6
+ bl_6 br_6 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_7
+ bl_7 br_7 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_8
+ bl_8 br_8 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_9
+ bl_9 br_9 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_10
+ bl_10 br_10 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_11
+ bl_11 br_11 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_12
+ bl_12 br_12 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_13
+ bl_13 br_13 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_14
+ bl_14 br_14 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_15
+ bl_15 br_15 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_16
+ bl_16 br_16 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_17
+ bl_17 br_17 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_18
+ bl_18 br_18 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_19
+ bl_19 br_19 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_20
+ bl_20 br_20 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_21
+ bl_21 br_21 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_22
+ bl_22 br_22 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_23
+ bl_23 br_23 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_24
+ bl_24 br_24 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_25
+ bl_25 br_25 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_26
+ bl_26 br_26 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_27
+ bl_27 br_27 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_28
+ bl_28 br_28 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_29
+ bl_29 br_29 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_30
+ bl_30 br_30 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_31
+ bl_31 br_31 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_32
+ bl_32 br_32 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_33
+ bl_33 br_33 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_34
+ bl_34 br_34 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_35
+ bl_35 br_35 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_36
+ bl_36 br_36 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_37
+ bl_37 br_37 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_38
+ bl_38 br_38 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_39
+ bl_39 br_39 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_40
+ bl_40 br_40 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_41
+ bl_41 br_41 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_42
+ bl_42 br_42 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_43
+ bl_43 br_43 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_44
+ bl_44 br_44 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_45
+ bl_45 br_45 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_46
+ bl_46 br_46 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_47
+ bl_47 br_47 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_48
+ bl_48 br_48 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_49
+ bl_49 br_49 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_50
+ bl_50 br_50 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_51
+ bl_51 br_51 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_52
+ bl_52 br_52 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_53
+ bl_53 br_53 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_54
+ bl_54 br_54 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_55
+ bl_55 br_55 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_56
+ bl_56 br_56 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_57
+ bl_57 br_57 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_58
+ bl_58 br_58 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_59
+ bl_59 br_59 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_60
+ bl_60 br_60 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_61
+ bl_61 br_61 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_62
+ bl_62 br_62 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_63
+ bl_63 br_63 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_64
+ bl_64 br_64 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_65
+ bl_65 br_65 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_66
+ bl_66 br_66 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_67
+ bl_67 br_67 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_68
+ bl_68 br_68 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_69
+ bl_69 br_69 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_70
+ bl_70 br_70 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_71
+ bl_71 br_71 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_72
+ bl_72 br_72 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_73
+ bl_73 br_73 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_74
+ bl_74 br_74 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_75
+ bl_75 br_75 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_76
+ bl_76 br_76 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_77
+ bl_77 br_77 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_78
+ bl_78 br_78 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_79
+ bl_79 br_79 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_80
+ bl_80 br_80 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_81
+ bl_81 br_81 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_82
+ bl_82 br_82 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_83
+ bl_83 br_83 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_84
+ bl_84 br_84 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_85
+ bl_85 br_85 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_86
+ bl_86 br_86 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_87
+ bl_87 br_87 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_88
+ bl_88 br_88 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_89
+ bl_89 br_89 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_90
+ bl_90 br_90 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_91
+ bl_91 br_91 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_92
+ bl_92 br_92 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_93
+ bl_93 br_93 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_94
+ bl_94 br_94 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_95
+ bl_95 br_95 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_96
+ bl_96 br_96 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_97
+ bl_97 br_97 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_98
+ bl_98 br_98 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_99
+ bl_99 br_99 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_100
+ bl_100 br_100 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_101
+ bl_101 br_101 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_102
+ bl_102 br_102 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_103
+ bl_103 br_103 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_104
+ bl_104 br_104 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_105
+ bl_105 br_105 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_106
+ bl_106 br_106 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_107
+ bl_107 br_107 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_108
+ bl_108 br_108 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_109
+ bl_109 br_109 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_110
+ bl_110 br_110 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_111
+ bl_111 br_111 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_112
+ bl_112 br_112 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_113
+ bl_113 br_113 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_114
+ bl_114 br_114 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_115
+ bl_115 br_115 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_116
+ bl_116 br_116 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_117
+ bl_117 br_117 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_118
+ bl_118 br_118 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_119
+ bl_119 br_119 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_120
+ bl_120 br_120 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_121
+ bl_121 br_121 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_122
+ bl_122 br_122 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_123
+ bl_123 br_123 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_124
+ bl_124 br_124 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_125
+ bl_125 br_125 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_126
+ bl_126 br_126 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_127
+ bl_127 br_127 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_128
+ bl_128 br_128 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
Xpre_column_129
+ bl_129 br_129 en_bar vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_0
.ENDS sky130_sram_1kbyte_1rw_32x256_8_precharge_array

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_port_data
+ rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5
+ br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11
+ bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22
+ bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28
+ br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33
+ bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39
+ br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44
+ bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50
+ br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55
+ bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61
+ br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66
+ bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72
+ br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77
+ bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83
+ br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88
+ bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94
+ br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99
+ bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104
+ bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109
+ bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114
+ bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119
+ bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124
+ bl_125 br_125 bl_126 br_126 bl_127 br_127 sparebl_0 sparebr_0 dout_0
+ dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10
+ dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18
+ dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26
+ dout_27 dout_28 dout_29 dout_30 dout_31 dout_32 din_0 din_1 din_2
+ din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13
+ din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23
+ din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 din_32 sel_0
+ sel_1 sel_2 sel_3 s_en p_en_bar w_en bank_wmask_0 bank_wmask_1
+ bank_wmask_2 bank_wmask_3 bank_spare_wen0 vdd gnd
* INOUT : rbl_bl 
* INOUT : rbl_br 
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : sparebl_0 
* INOUT : sparebr_0 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* OUTPUT: dout_32 
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : din_32 
* INPUT : sel_0 
* INPUT : sel_1 
* INPUT : sel_2 
* INPUT : sel_3 
* INPUT : s_en 
* INPUT : p_en_bar 
* INPUT : w_en 
* INPUT : bank_wmask_0 
* INPUT : bank_wmask_1 
* INPUT : bank_wmask_2 
* INPUT : bank_wmask_3 
* INPUT : bank_spare_wen0 
* POWER : vdd 
* GROUND: gnd 
Xprecharge_array0
+ rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5
+ br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11
+ bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22
+ bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28
+ br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33
+ bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39
+ br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44
+ bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50
+ br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55
+ bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61
+ br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66
+ bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72
+ br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77
+ bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83
+ br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88
+ bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94
+ br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99
+ bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104
+ bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109
+ bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114
+ bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119
+ bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124
+ bl_125 br_125 bl_126 br_126 bl_127 br_127 sparebl_0 sparebr_0 p_en_bar
+ vdd
+ sky130_sram_1kbyte_1rw_32x256_8_precharge_array
Xsense_amp_array0
+ dout_0 bl_out_0 br_out_0 dout_1 bl_out_1 br_out_1 dout_2 bl_out_2
+ br_out_2 dout_3 bl_out_3 br_out_3 dout_4 bl_out_4 br_out_4 dout_5
+ bl_out_5 br_out_5 dout_6 bl_out_6 br_out_6 dout_7 bl_out_7 br_out_7
+ dout_8 bl_out_8 br_out_8 dout_9 bl_out_9 br_out_9 dout_10 bl_out_10
+ br_out_10 dout_11 bl_out_11 br_out_11 dout_12 bl_out_12 br_out_12
+ dout_13 bl_out_13 br_out_13 dout_14 bl_out_14 br_out_14 dout_15
+ bl_out_15 br_out_15 dout_16 bl_out_16 br_out_16 dout_17 bl_out_17
+ br_out_17 dout_18 bl_out_18 br_out_18 dout_19 bl_out_19 br_out_19
+ dout_20 bl_out_20 br_out_20 dout_21 bl_out_21 br_out_21 dout_22
+ bl_out_22 br_out_22 dout_23 bl_out_23 br_out_23 dout_24 bl_out_24
+ br_out_24 dout_25 bl_out_25 br_out_25 dout_26 bl_out_26 br_out_26
+ dout_27 bl_out_27 br_out_27 dout_28 bl_out_28 br_out_28 dout_29
+ bl_out_29 br_out_29 dout_30 bl_out_30 br_out_30 dout_31 bl_out_31
+ br_out_31 dout_32 sparebl_0 sparebr_0 s_en vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_sense_amp_array
Xwrite_driver_array0
+ din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10
+ din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20
+ din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30
+ din_31 din_32 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2
+ bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6
+ br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9
+ bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13
+ br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16
+ bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20
+ br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23
+ bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27
+ br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30
+ bl_out_31 br_out_31 sparebl_0 sparebr_0 wdriver_sel_0 wdriver_sel_1
+ wdriver_sel_2 wdriver_sel_3 bank_spare_wen0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_write_driver_array
Xwrite_mask_and_array0
+ bank_wmask_0 bank_wmask_1 bank_wmask_2 bank_wmask_3 w_en wdriver_sel_0
+ wdriver_sel_1 wdriver_sel_2 wdriver_sel_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_write_mask_and_array
Xcolumn_mux_array0
+ bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18
+ br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23
+ bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34
+ bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40
+ br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51
+ br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67
+ bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73
+ br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78
+ bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84
+ br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89
+ bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95
+ br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100
+ bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105
+ bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110
+ bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115
+ bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120
+ bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125
+ bl_126 br_126 bl_127 br_127 sel_0 sel_1 sel_2 sel_3 bl_out_0 br_out_0
+ bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4
+ br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7
+ bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11
+ br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14
+ bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18
+ br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21
+ bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25
+ br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28
+ bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_mux_array
.ENDS sky130_sram_1kbyte_1rw_32x256_8_port_data

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_dec_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 32
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_dec_0
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* NGSPICE file created from sky130_fd_bd_sram__openram_sp_nand2_dec.ext - technology: EFS8A


* Top level circuit sky130_fd_bd_sram__openram_sp_nand2_dec
.subckt sky130_fd_bd_sram__openram_sp_nand2_dec A B Z VDD GND

X1001 Z B VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1002 VDD A Z VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1000 Z A a_n722_276# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1003 a_n722_276# B GND GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
.ends


.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* cols: 129
Xwld_nand
+ A B zb_int vdd gnd
+ sky130_fd_bd_sram__openram_sp_nand2_dec
Xwl_driver
+ zb_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_dec_0
.ENDS sky130_sram_1kbyte_1rw_32x256_8_wordline_driver

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_wordline_driver_array
+ in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12
+ in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23
+ in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34
+ in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45
+ in_46 in_47 in_48 in_49 in_50 in_51 in_52 in_53 in_54 in_55 in_56
+ in_57 in_58 in_59 in_60 in_61 in_62 in_63 in_64 wl_0 wl_1 wl_2 wl_3
+ wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26
+ wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37
+ wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48
+ wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59
+ wl_60 wl_61 wl_62 wl_63 wl_64 en vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* INPUT : in_32 
* INPUT : in_33 
* INPUT : in_34 
* INPUT : in_35 
* INPUT : in_36 
* INPUT : in_37 
* INPUT : in_38 
* INPUT : in_39 
* INPUT : in_40 
* INPUT : in_41 
* INPUT : in_42 
* INPUT : in_43 
* INPUT : in_44 
* INPUT : in_45 
* INPUT : in_46 
* INPUT : in_47 
* INPUT : in_48 
* INPUT : in_49 
* INPUT : in_50 
* INPUT : in_51 
* INPUT : in_52 
* INPUT : in_53 
* INPUT : in_54 
* INPUT : in_55 
* INPUT : in_56 
* INPUT : in_57 
* INPUT : in_58 
* INPUT : in_59 
* INPUT : in_60 
* INPUT : in_61 
* INPUT : in_62 
* INPUT : in_63 
* INPUT : in_64 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* rows: 65 cols: 129
Xwl_driver_and0
+ in_0 en wl_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and1
+ in_1 en wl_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and2
+ in_2 en wl_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and3
+ in_3 en wl_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and4
+ in_4 en wl_4 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and5
+ in_5 en wl_5 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and6
+ in_6 en wl_6 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and7
+ in_7 en wl_7 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and8
+ in_8 en wl_8 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and9
+ in_9 en wl_9 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and10
+ in_10 en wl_10 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and11
+ in_11 en wl_11 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and12
+ in_12 en wl_12 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and13
+ in_13 en wl_13 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and14
+ in_14 en wl_14 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and15
+ in_15 en wl_15 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and16
+ in_16 en wl_16 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and17
+ in_17 en wl_17 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and18
+ in_18 en wl_18 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and19
+ in_19 en wl_19 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and20
+ in_20 en wl_20 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and21
+ in_21 en wl_21 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and22
+ in_22 en wl_22 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and23
+ in_23 en wl_23 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and24
+ in_24 en wl_24 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and25
+ in_25 en wl_25 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and26
+ in_26 en wl_26 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and27
+ in_27 en wl_27 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and28
+ in_28 en wl_28 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and29
+ in_29 en wl_29 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and30
+ in_30 en wl_30 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and31
+ in_31 en wl_31 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and32
+ in_32 en wl_32 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and33
+ in_33 en wl_33 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and34
+ in_34 en wl_34 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and35
+ in_35 en wl_35 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and36
+ in_36 en wl_36 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and37
+ in_37 en wl_37 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and38
+ in_38 en wl_38 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and39
+ in_39 en wl_39 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and40
+ in_40 en wl_40 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and41
+ in_41 en wl_41 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and42
+ in_42 en wl_42 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and43
+ in_43 en wl_43 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and44
+ in_44 en wl_44 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and45
+ in_45 en wl_45 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and46
+ in_46 en wl_46 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and47
+ in_47 en wl_47 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and48
+ in_48 en wl_48 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and49
+ in_49 en wl_49 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and50
+ in_50 en wl_50 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and51
+ in_51 en wl_51 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and52
+ in_52 en wl_52 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and53
+ in_53 en wl_53 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and54
+ in_54 en wl_54 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and55
+ in_55 en wl_55 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and56
+ in_56 en wl_56 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and57
+ in_57 en wl_57 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and58
+ in_58 en wl_58 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and59
+ in_59 en wl_59 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and60
+ in_60 en wl_60 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and61
+ in_61 en wl_61 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and62
+ in_62 en wl_62 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and63
+ in_63 en wl_63 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
Xwl_driver_and64
+ in_64 en wl_64 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver
.ENDS sky130_sram_1kbyte_1rw_32x256_8_wordline_driver_array

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_and2_dec_0
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 32
Xpand2_dec_nand
+ A B zb_int vdd gnd
+ sky130_fd_bd_sram__openram_sp_nand2_dec
Xpand2_dec_inv
+ zb_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_dec_0
.ENDS sky130_sram_1kbyte_1rw_32x256_8_and2_dec_0

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_pinv_dec
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS sky130_sram_1kbyte_1rw_32x256_8_pinv_dec

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_and2_dec
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand2_dec_nand
+ A B zb_int vdd gnd
+ sky130_fd_bd_sram__openram_sp_nand2_dec
Xpand2_dec_inv
+ zb_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_dec
.ENDS sky130_sram_1kbyte_1rw_32x256_8_and2_dec

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_hierarchical_predecode2x4
+ in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0
+ in_0 inbar_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_dec
Xpre_inv_1
+ in_1 inbar_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_dec
XXpre2x4_and_0
+ inbar_0 inbar_1 out_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and2_dec
XXpre2x4_and_1
+ in_0 inbar_1 out_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and2_dec
XXpre2x4_and_2
+ inbar_0 in_1 out_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and2_dec
XXpre2x4_and_3
+ in_0 in_1 out_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and2_dec
.ENDS sky130_sram_1kbyte_1rw_32x256_8_hierarchical_predecode2x4
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* NGSPICE file created from sky130_fd_bd_sram__openram_sp_nand3_dec.ext - technology: EFS8A


* Top level circuit sky130_fd_bd_sram__openram_sp_nand3_dec
.subckt sky130_fd_bd_sram__openram_sp_nand3_dec A B C Z VDD GND

X1001 Z A a_n346_328# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1002 a_n346_256# C GND GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1003 a_n346_328# B a_n346_256# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1000 Z B VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1004 Z A VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1005 Z C VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
.ends


.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_and3_dec
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand3_dec_nand
+ A B C zb_int vdd gnd
+ sky130_fd_bd_sram__openram_sp_nand3_dec
Xpand3_dec_inv
+ zb_int Z vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_dec
.ENDS sky130_sram_1kbyte_1rw_32x256_8_and3_dec

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_hierarchical_predecode3x8
+ in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0
+ in_0 inbar_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_dec
Xpre_inv_1
+ in_1 inbar_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_dec
Xpre_inv_2
+ in_2 inbar_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_pinv_dec
XXpre3x8_and_0
+ inbar_0 inbar_1 inbar_2 out_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XXpre3x8_and_1
+ in_0 inbar_1 inbar_2 out_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XXpre3x8_and_2
+ inbar_0 in_1 inbar_2 out_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XXpre3x8_and_3
+ in_0 in_1 inbar_2 out_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XXpre3x8_and_4
+ inbar_0 inbar_1 in_2 out_4 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XXpre3x8_and_5
+ in_0 inbar_1 in_2 out_5 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XXpre3x8_and_6
+ inbar_0 in_1 in_2 out_6 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XXpre3x8_and_7
+ in_0 in_1 in_2 out_7 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
.ENDS sky130_sram_1kbyte_1rw_32x256_8_hierarchical_predecode3x8

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_hierarchical_decoder
+ addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 decode_0 decode_1
+ decode_2 decode_3 decode_4 decode_5 decode_6 decode_7 decode_8
+ decode_9 decode_10 decode_11 decode_12 decode_13 decode_14 decode_15
+ decode_16 decode_17 decode_18 decode_19 decode_20 decode_21 decode_22
+ decode_23 decode_24 decode_25 decode_26 decode_27 decode_28 decode_29
+ decode_30 decode_31 decode_32 decode_33 decode_34 decode_35 decode_36
+ decode_37 decode_38 decode_39 decode_40 decode_41 decode_42 decode_43
+ decode_44 decode_45 decode_46 decode_47 decode_48 decode_49 decode_50
+ decode_51 decode_52 decode_53 decode_54 decode_55 decode_56 decode_57
+ decode_58 decode_59 decode_60 decode_61 decode_62 decode_63 decode_64
+ vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* OUTPUT: decode_0 
* OUTPUT: decode_1 
* OUTPUT: decode_2 
* OUTPUT: decode_3 
* OUTPUT: decode_4 
* OUTPUT: decode_5 
* OUTPUT: decode_6 
* OUTPUT: decode_7 
* OUTPUT: decode_8 
* OUTPUT: decode_9 
* OUTPUT: decode_10 
* OUTPUT: decode_11 
* OUTPUT: decode_12 
* OUTPUT: decode_13 
* OUTPUT: decode_14 
* OUTPUT: decode_15 
* OUTPUT: decode_16 
* OUTPUT: decode_17 
* OUTPUT: decode_18 
* OUTPUT: decode_19 
* OUTPUT: decode_20 
* OUTPUT: decode_21 
* OUTPUT: decode_22 
* OUTPUT: decode_23 
* OUTPUT: decode_24 
* OUTPUT: decode_25 
* OUTPUT: decode_26 
* OUTPUT: decode_27 
* OUTPUT: decode_28 
* OUTPUT: decode_29 
* OUTPUT: decode_30 
* OUTPUT: decode_31 
* OUTPUT: decode_32 
* OUTPUT: decode_33 
* OUTPUT: decode_34 
* OUTPUT: decode_35 
* OUTPUT: decode_36 
* OUTPUT: decode_37 
* OUTPUT: decode_38 
* OUTPUT: decode_39 
* OUTPUT: decode_40 
* OUTPUT: decode_41 
* OUTPUT: decode_42 
* OUTPUT: decode_43 
* OUTPUT: decode_44 
* OUTPUT: decode_45 
* OUTPUT: decode_46 
* OUTPUT: decode_47 
* OUTPUT: decode_48 
* OUTPUT: decode_49 
* OUTPUT: decode_50 
* OUTPUT: decode_51 
* OUTPUT: decode_52 
* OUTPUT: decode_53 
* OUTPUT: decode_54 
* OUTPUT: decode_55 
* OUTPUT: decode_56 
* OUTPUT: decode_57 
* OUTPUT: decode_58 
* OUTPUT: decode_59 
* OUTPUT: decode_60 
* OUTPUT: decode_61 
* OUTPUT: decode_62 
* OUTPUT: decode_63 
* OUTPUT: decode_64 
* POWER : vdd 
* GROUND: gnd 
Xpre_0
+ addr_0 addr_1 out_0 out_1 out_2 out_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_hierarchical_predecode2x4
Xpre_1
+ addr_2 addr_3 out_4 out_5 out_6 out_7 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_hierarchical_predecode2x4
Xpre3x8_0
+ addr_4 addr_5 addr_6 out_8 out_9 out_10 out_11 out_12 out_13 out_14
+ out_15 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_hierarchical_predecode3x8
XDEC_AND_0
+ out_0 out_4 out_8 decode_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_16
+ out_0 out_4 out_9 decode_16 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_32
+ out_0 out_4 out_10 decode_32 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_48
+ out_0 out_4 out_11 decode_48 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_64
+ out_0 out_4 out_12 decode_64 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_4
+ out_0 out_5 out_8 decode_4 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_20
+ out_0 out_5 out_9 decode_20 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_36
+ out_0 out_5 out_10 decode_36 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_52
+ out_0 out_5 out_11 decode_52 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_8
+ out_0 out_6 out_8 decode_8 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_24
+ out_0 out_6 out_9 decode_24 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_40
+ out_0 out_6 out_10 decode_40 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_56
+ out_0 out_6 out_11 decode_56 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_12
+ out_0 out_7 out_8 decode_12 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_28
+ out_0 out_7 out_9 decode_28 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_44
+ out_0 out_7 out_10 decode_44 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_60
+ out_0 out_7 out_11 decode_60 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_1
+ out_1 out_4 out_8 decode_1 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_17
+ out_1 out_4 out_9 decode_17 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_33
+ out_1 out_4 out_10 decode_33 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_49
+ out_1 out_4 out_11 decode_49 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_5
+ out_1 out_5 out_8 decode_5 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_21
+ out_1 out_5 out_9 decode_21 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_37
+ out_1 out_5 out_10 decode_37 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_53
+ out_1 out_5 out_11 decode_53 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_9
+ out_1 out_6 out_8 decode_9 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_25
+ out_1 out_6 out_9 decode_25 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_41
+ out_1 out_6 out_10 decode_41 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_57
+ out_1 out_6 out_11 decode_57 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_13
+ out_1 out_7 out_8 decode_13 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_29
+ out_1 out_7 out_9 decode_29 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_45
+ out_1 out_7 out_10 decode_45 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_61
+ out_1 out_7 out_11 decode_61 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_2
+ out_2 out_4 out_8 decode_2 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_18
+ out_2 out_4 out_9 decode_18 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_34
+ out_2 out_4 out_10 decode_34 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_50
+ out_2 out_4 out_11 decode_50 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_6
+ out_2 out_5 out_8 decode_6 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_22
+ out_2 out_5 out_9 decode_22 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_38
+ out_2 out_5 out_10 decode_38 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_54
+ out_2 out_5 out_11 decode_54 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_10
+ out_2 out_6 out_8 decode_10 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_26
+ out_2 out_6 out_9 decode_26 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_42
+ out_2 out_6 out_10 decode_42 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_58
+ out_2 out_6 out_11 decode_58 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_14
+ out_2 out_7 out_8 decode_14 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_30
+ out_2 out_7 out_9 decode_30 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_46
+ out_2 out_7 out_10 decode_46 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_62
+ out_2 out_7 out_11 decode_62 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_3
+ out_3 out_4 out_8 decode_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_19
+ out_3 out_4 out_9 decode_19 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_35
+ out_3 out_4 out_10 decode_35 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_51
+ out_3 out_4 out_11 decode_51 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_7
+ out_3 out_5 out_8 decode_7 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_23
+ out_3 out_5 out_9 decode_23 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_39
+ out_3 out_5 out_10 decode_39 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_55
+ out_3 out_5 out_11 decode_55 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_11
+ out_3 out_6 out_8 decode_11 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_27
+ out_3 out_6 out_9 decode_27 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_43
+ out_3 out_6 out_10 decode_43 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_59
+ out_3 out_6 out_11 decode_59 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_15
+ out_3 out_7 out_8 decode_15 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_31
+ out_3 out_7 out_9 decode_31 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_47
+ out_3 out_7 out_10 decode_47 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
XDEC_AND_63
+ out_3 out_7 out_11 decode_63 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and3_dec
.ENDS sky130_sram_1kbyte_1rw_32x256_8_hierarchical_decoder

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_port_address
+ addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 wl_en wl_0 wl_1 wl_2
+ wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26
+ wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37
+ wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48
+ wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59
+ wl_60 wl_61 wl_62 wl_63 wl_64 rbl_wl vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* INPUT : wl_en 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: rbl_wl 
* POWER : vdd 
* GROUND: gnd 
Xrow_decoder
+ addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 dec_out_0 dec_out_1
+ dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8
+ dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14
+ dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20
+ dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26
+ dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32
+ dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38
+ dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44
+ dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50
+ dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56
+ dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62
+ dec_out_63 dec_out_64 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_hierarchical_decoder
Xwordline_driver
+ dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6
+ dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12
+ dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18
+ dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24
+ dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30
+ dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36
+ dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42
+ dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48
+ dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54
+ dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60
+ dec_out_61 dec_out_62 dec_out_63 dec_out_64 wl_0 wl_1 wl_2 wl_3 wl_4
+ wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16
+ wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27
+ wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38
+ wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49
+ wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60
+ wl_61 wl_62 wl_63 wl_64 wl_en vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_wordline_driver_array
Xrbl_driver
+ wl_en vdd rbl_wl vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_and2_dec_0
.ENDS sky130_sram_1kbyte_1rw_32x256_8_port_address
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_wlstrap_p.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_wlstrap_p VGND
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_wlstrapa_p.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_wlstrapa_p VGND
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colend.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colend bl vdd gnd br gate vpb vnb
*X0 br gate br vnb sky130_fd_pr__special_nfet_pass w=0.07u l=0.21u
.ends

* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colend_p_cent.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colend_p_cent VGND VPB VNB
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colenda.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colenda bl vdd gnd br gate vpb vnb
*X0 br gate br vnb sky130_fd_pr__special_nfet_pass w=0.065u l=0.17u
.ends

* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_opt1a_replica.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_cell_opt1a_replica BL BR VGND VPWR VPB VNB WL
X0 VPWR WL BR VNB sky130_fd_pr__special_nfet_pass ad=4.375e+10p pd=920000u as=1.68e+10p ps=520000u w=140000u l=150000u
X1 Q VPWR VGND VNB sky130_fd_pr__special_nfet_latch ad=1.56e+11p pd=2.38e+06u as=8.08e+10p ps=1.28e+06u w=210000u l=150000u
X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass ad=1.68e+10p pd=520000u as=4.25e+10p ps=920000u w=140000u l=150000u
*X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass ad=3.5e+10p pd=780000u as=0p ps=0u w=70000u l=95000u
*X4 VPWR WL VPWR VPB sky130_fd_pr__special_pfet_pass ad=9.72e+10p pd=1.86e+06u as=0p ps=0u w=70000u l=95000u
X5 VPWR Q VPWR VPB sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X6 Q VPWR VPWR VPB sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X7 VGND Q VPWR VNB sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colenda_p_cent.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colenda_p_cent VGND VPB VNB
.ends
* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_opt1_replica.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_cell_opt1_replica BL BR VGND VPWR VPB VNB WL
X0 VPWR WL BR VNB sky130_fd_pr__special_nfet_pass ad=4.375e+10p pd=920000u as=1.68e+10p ps=520000u w=140000u l=150000u
X1 Q VPWR VGND VNB sky130_fd_pr__special_nfet_latch ad=1.56e+11p pd=2.38e+06u as=8.08e+10p ps=1.28e+06u w=210000u l=150000u
X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass ad=1.68e+10p pd=520000u as=4.25e+10p ps=920000u w=140000u l=150000u
*X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass ad=3.5e+10p pd=780000u as=0p ps=0u w=70000u l=95000u
*X4 VPWR WL VPWR VPB sky130_fd_pr__special_pfet_pass ad=9.72e+10p pd=1.86e+06u as=0p ps=0u w=70000u l=95000u
X5 VPWR Q VPWR VPB sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X6 Q VPWR VPWR VPB sky130_fd_pr__special_pfet_pass ad=0p pd=0u as=0p ps=0u w=140000u l=150000u
X7 VGND Q VPWR VNB sky130_fd_pr__special_nfet_latch ad=0p pd=0u as=0p ps=0u w=210000u l=150000u
.ends

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_sky130_replica_column
+ bl_0_0 br_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8
+ wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17
+ wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25
+ wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33
+ wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41
+ wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49
+ wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57
+ wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65
+ wl_0_66 vdd gnd top_gate bot_gate
* OUTPUT: bl_0_0 
* OUTPUT: br_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* POWER : vdd 
* GROUND: gnd 
* INPUT : top_gate 
* INPUT : bot_gate 
Xrbc_0
+ bl_0_0 vdd gnd br_0_0 top_gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrbc_0_cap
+ gnd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrbc_1
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_1_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_2
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_2_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_3
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_3_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_4
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_4_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_5
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_5_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_6
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_6_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_7
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_7_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_8
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_8_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_9
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_9_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_10
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_10_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_11
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_11_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_12
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_12_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_13
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_13_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_14
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_14_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_15
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_15_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_16
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_16_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_17
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_17_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_18
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_18_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_19
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_19_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_20
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_20_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_21
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_21_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_22
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_22_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_23
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_23_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_24
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_24_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_25
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_25_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_26
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_26_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_27
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_27_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_28
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_28_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_29
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_29_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_30
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_30_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_31
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_31_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_32
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_32_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_33
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_33_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_34
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_34_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_35
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_35_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_36
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_36_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_37
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_37_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_38
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_38_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_39
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_39_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_40
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_40_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_41
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_41_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_42
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_42_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_43
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_43_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_44
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_44_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_45
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_45_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_46
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_46_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_47
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_47_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_48
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_48_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_49
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_49_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_50
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_50_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_51
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_51_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_52
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_52_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_53
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_53_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_54
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_54_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_55
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_55_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_56
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_56_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_57
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_57_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_58
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_58_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_59
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_59_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_60
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_60_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_61
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_61_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_62
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_62_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_63
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_63_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_64
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_64_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_65
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_65
+ sky130_fd_bd_sram__openram_sp_cell_opt1_replica
Xrbc_65_strap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrbc_66
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_66
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_replica
Xrbc_66_strap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrbc_67
+ bl_0_0 vdd gnd br_0_0 bot_gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrbc_67_cap
+ gnd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
.ENDS sky130_sram_1kbyte_1rw_32x256_8_sky130_replica_column
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colenda_cent.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colenda_cent VPWR VPB VNB
.ends

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_sky130_col_cap_array_0
+ fake_bl_0 fake_br_0 fake_bl_1 fake_br_1 fake_bl_2 fake_br_2 fake_bl_3
+ fake_br_3 fake_bl_4 fake_br_4 fake_bl_5 fake_br_5 fake_bl_6 fake_br_6
+ fake_bl_7 fake_br_7 fake_bl_8 fake_br_8 fake_bl_9 fake_br_9 fake_bl_10
+ fake_br_10 fake_bl_11 fake_br_11 fake_bl_12 fake_br_12 fake_bl_13
+ fake_br_13 fake_bl_14 fake_br_14 fake_bl_15 fake_br_15 fake_bl_16
+ fake_br_16 fake_bl_17 fake_br_17 fake_bl_18 fake_br_18 fake_bl_19
+ fake_br_19 fake_bl_20 fake_br_20 fake_bl_21 fake_br_21 fake_bl_22
+ fake_br_22 fake_bl_23 fake_br_23 fake_bl_24 fake_br_24 fake_bl_25
+ fake_br_25 fake_bl_26 fake_br_26 fake_bl_27 fake_br_27 fake_bl_28
+ fake_br_28 fake_bl_29 fake_br_29 fake_bl_30 fake_br_30 fake_bl_31
+ fake_br_31 fake_bl_32 fake_br_32 fake_bl_33 fake_br_33 fake_bl_34
+ fake_br_34 fake_bl_35 fake_br_35 fake_bl_36 fake_br_36 fake_bl_37
+ fake_br_37 fake_bl_38 fake_br_38 fake_bl_39 fake_br_39 fake_bl_40
+ fake_br_40 fake_bl_41 fake_br_41 fake_bl_42 fake_br_42 fake_bl_43
+ fake_br_43 fake_bl_44 fake_br_44 fake_bl_45 fake_br_45 fake_bl_46
+ fake_br_46 fake_bl_47 fake_br_47 fake_bl_48 fake_br_48 fake_bl_49
+ fake_br_49 fake_bl_50 fake_br_50 fake_bl_51 fake_br_51 fake_bl_52
+ fake_br_52 fake_bl_53 fake_br_53 fake_bl_54 fake_br_54 fake_bl_55
+ fake_br_55 fake_bl_56 fake_br_56 fake_bl_57 fake_br_57 fake_bl_58
+ fake_br_58 fake_bl_59 fake_br_59 fake_bl_60 fake_br_60 fake_bl_61
+ fake_br_61 fake_bl_62 fake_br_62 fake_bl_63 fake_br_63 fake_bl_64
+ fake_br_64 fake_bl_65 fake_br_65 fake_bl_66 fake_br_66 fake_bl_67
+ fake_br_67 fake_bl_68 fake_br_68 fake_bl_69 fake_br_69 fake_bl_70
+ fake_br_70 fake_bl_71 fake_br_71 fake_bl_72 fake_br_72 fake_bl_73
+ fake_br_73 fake_bl_74 fake_br_74 fake_bl_75 fake_br_75 fake_bl_76
+ fake_br_76 fake_bl_77 fake_br_77 fake_bl_78 fake_br_78 fake_bl_79
+ fake_br_79 fake_bl_80 fake_br_80 fake_bl_81 fake_br_81 fake_bl_82
+ fake_br_82 fake_bl_83 fake_br_83 fake_bl_84 fake_br_84 fake_bl_85
+ fake_br_85 fake_bl_86 fake_br_86 fake_bl_87 fake_br_87 fake_bl_88
+ fake_br_88 fake_bl_89 fake_br_89 fake_bl_90 fake_br_90 fake_bl_91
+ fake_br_91 fake_bl_92 fake_br_92 fake_bl_93 fake_br_93 fake_bl_94
+ fake_br_94 fake_bl_95 fake_br_95 fake_bl_96 fake_br_96 fake_bl_97
+ fake_br_97 fake_bl_98 fake_br_98 fake_bl_99 fake_br_99 fake_bl_100
+ fake_br_100 fake_bl_101 fake_br_101 fake_bl_102 fake_br_102
+ fake_bl_103 fake_br_103 fake_bl_104 fake_br_104 fake_bl_105
+ fake_br_105 fake_bl_106 fake_br_106 fake_bl_107 fake_br_107
+ fake_bl_108 fake_br_108 fake_bl_109 fake_br_109 fake_bl_110
+ fake_br_110 fake_bl_111 fake_br_111 fake_bl_112 fake_br_112
+ fake_bl_113 fake_br_113 fake_bl_114 fake_br_114 fake_bl_115
+ fake_br_115 fake_bl_116 fake_br_116 fake_bl_117 fake_br_117
+ fake_bl_118 fake_br_118 fake_bl_119 fake_br_119 fake_bl_120
+ fake_br_120 fake_bl_121 fake_br_121 fake_bl_122 fake_br_122
+ fake_bl_123 fake_br_123 fake_bl_124 fake_br_124 fake_bl_125
+ fake_br_125 fake_bl_126 fake_br_126 fake_bl_127 fake_br_127
+ fake_bl_128 fake_br_128 vdd gnd gate
* OUTPUT: fake_bl_0 
* OUTPUT: fake_br_0 
* OUTPUT: fake_bl_1 
* OUTPUT: fake_br_1 
* OUTPUT: fake_bl_2 
* OUTPUT: fake_br_2 
* OUTPUT: fake_bl_3 
* OUTPUT: fake_br_3 
* OUTPUT: fake_bl_4 
* OUTPUT: fake_br_4 
* OUTPUT: fake_bl_5 
* OUTPUT: fake_br_5 
* OUTPUT: fake_bl_6 
* OUTPUT: fake_br_6 
* OUTPUT: fake_bl_7 
* OUTPUT: fake_br_7 
* OUTPUT: fake_bl_8 
* OUTPUT: fake_br_8 
* OUTPUT: fake_bl_9 
* OUTPUT: fake_br_9 
* OUTPUT: fake_bl_10 
* OUTPUT: fake_br_10 
* OUTPUT: fake_bl_11 
* OUTPUT: fake_br_11 
* OUTPUT: fake_bl_12 
* OUTPUT: fake_br_12 
* OUTPUT: fake_bl_13 
* OUTPUT: fake_br_13 
* OUTPUT: fake_bl_14 
* OUTPUT: fake_br_14 
* OUTPUT: fake_bl_15 
* OUTPUT: fake_br_15 
* OUTPUT: fake_bl_16 
* OUTPUT: fake_br_16 
* OUTPUT: fake_bl_17 
* OUTPUT: fake_br_17 
* OUTPUT: fake_bl_18 
* OUTPUT: fake_br_18 
* OUTPUT: fake_bl_19 
* OUTPUT: fake_br_19 
* OUTPUT: fake_bl_20 
* OUTPUT: fake_br_20 
* OUTPUT: fake_bl_21 
* OUTPUT: fake_br_21 
* OUTPUT: fake_bl_22 
* OUTPUT: fake_br_22 
* OUTPUT: fake_bl_23 
* OUTPUT: fake_br_23 
* OUTPUT: fake_bl_24 
* OUTPUT: fake_br_24 
* OUTPUT: fake_bl_25 
* OUTPUT: fake_br_25 
* OUTPUT: fake_bl_26 
* OUTPUT: fake_br_26 
* OUTPUT: fake_bl_27 
* OUTPUT: fake_br_27 
* OUTPUT: fake_bl_28 
* OUTPUT: fake_br_28 
* OUTPUT: fake_bl_29 
* OUTPUT: fake_br_29 
* OUTPUT: fake_bl_30 
* OUTPUT: fake_br_30 
* OUTPUT: fake_bl_31 
* OUTPUT: fake_br_31 
* OUTPUT: fake_bl_32 
* OUTPUT: fake_br_32 
* OUTPUT: fake_bl_33 
* OUTPUT: fake_br_33 
* OUTPUT: fake_bl_34 
* OUTPUT: fake_br_34 
* OUTPUT: fake_bl_35 
* OUTPUT: fake_br_35 
* OUTPUT: fake_bl_36 
* OUTPUT: fake_br_36 
* OUTPUT: fake_bl_37 
* OUTPUT: fake_br_37 
* OUTPUT: fake_bl_38 
* OUTPUT: fake_br_38 
* OUTPUT: fake_bl_39 
* OUTPUT: fake_br_39 
* OUTPUT: fake_bl_40 
* OUTPUT: fake_br_40 
* OUTPUT: fake_bl_41 
* OUTPUT: fake_br_41 
* OUTPUT: fake_bl_42 
* OUTPUT: fake_br_42 
* OUTPUT: fake_bl_43 
* OUTPUT: fake_br_43 
* OUTPUT: fake_bl_44 
* OUTPUT: fake_br_44 
* OUTPUT: fake_bl_45 
* OUTPUT: fake_br_45 
* OUTPUT: fake_bl_46 
* OUTPUT: fake_br_46 
* OUTPUT: fake_bl_47 
* OUTPUT: fake_br_47 
* OUTPUT: fake_bl_48 
* OUTPUT: fake_br_48 
* OUTPUT: fake_bl_49 
* OUTPUT: fake_br_49 
* OUTPUT: fake_bl_50 
* OUTPUT: fake_br_50 
* OUTPUT: fake_bl_51 
* OUTPUT: fake_br_51 
* OUTPUT: fake_bl_52 
* OUTPUT: fake_br_52 
* OUTPUT: fake_bl_53 
* OUTPUT: fake_br_53 
* OUTPUT: fake_bl_54 
* OUTPUT: fake_br_54 
* OUTPUT: fake_bl_55 
* OUTPUT: fake_br_55 
* OUTPUT: fake_bl_56 
* OUTPUT: fake_br_56 
* OUTPUT: fake_bl_57 
* OUTPUT: fake_br_57 
* OUTPUT: fake_bl_58 
* OUTPUT: fake_br_58 
* OUTPUT: fake_bl_59 
* OUTPUT: fake_br_59 
* OUTPUT: fake_bl_60 
* OUTPUT: fake_br_60 
* OUTPUT: fake_bl_61 
* OUTPUT: fake_br_61 
* OUTPUT: fake_bl_62 
* OUTPUT: fake_br_62 
* OUTPUT: fake_bl_63 
* OUTPUT: fake_br_63 
* OUTPUT: fake_bl_64 
* OUTPUT: fake_br_64 
* OUTPUT: fake_bl_65 
* OUTPUT: fake_br_65 
* OUTPUT: fake_bl_66 
* OUTPUT: fake_br_66 
* OUTPUT: fake_bl_67 
* OUTPUT: fake_br_67 
* OUTPUT: fake_bl_68 
* OUTPUT: fake_br_68 
* OUTPUT: fake_bl_69 
* OUTPUT: fake_br_69 
* OUTPUT: fake_bl_70 
* OUTPUT: fake_br_70 
* OUTPUT: fake_bl_71 
* OUTPUT: fake_br_71 
* OUTPUT: fake_bl_72 
* OUTPUT: fake_br_72 
* OUTPUT: fake_bl_73 
* OUTPUT: fake_br_73 
* OUTPUT: fake_bl_74 
* OUTPUT: fake_br_74 
* OUTPUT: fake_bl_75 
* OUTPUT: fake_br_75 
* OUTPUT: fake_bl_76 
* OUTPUT: fake_br_76 
* OUTPUT: fake_bl_77 
* OUTPUT: fake_br_77 
* OUTPUT: fake_bl_78 
* OUTPUT: fake_br_78 
* OUTPUT: fake_bl_79 
* OUTPUT: fake_br_79 
* OUTPUT: fake_bl_80 
* OUTPUT: fake_br_80 
* OUTPUT: fake_bl_81 
* OUTPUT: fake_br_81 
* OUTPUT: fake_bl_82 
* OUTPUT: fake_br_82 
* OUTPUT: fake_bl_83 
* OUTPUT: fake_br_83 
* OUTPUT: fake_bl_84 
* OUTPUT: fake_br_84 
* OUTPUT: fake_bl_85 
* OUTPUT: fake_br_85 
* OUTPUT: fake_bl_86 
* OUTPUT: fake_br_86 
* OUTPUT: fake_bl_87 
* OUTPUT: fake_br_87 
* OUTPUT: fake_bl_88 
* OUTPUT: fake_br_88 
* OUTPUT: fake_bl_89 
* OUTPUT: fake_br_89 
* OUTPUT: fake_bl_90 
* OUTPUT: fake_br_90 
* OUTPUT: fake_bl_91 
* OUTPUT: fake_br_91 
* OUTPUT: fake_bl_92 
* OUTPUT: fake_br_92 
* OUTPUT: fake_bl_93 
* OUTPUT: fake_br_93 
* OUTPUT: fake_bl_94 
* OUTPUT: fake_br_94 
* OUTPUT: fake_bl_95 
* OUTPUT: fake_br_95 
* OUTPUT: fake_bl_96 
* OUTPUT: fake_br_96 
* OUTPUT: fake_bl_97 
* OUTPUT: fake_br_97 
* OUTPUT: fake_bl_98 
* OUTPUT: fake_br_98 
* OUTPUT: fake_bl_99 
* OUTPUT: fake_br_99 
* OUTPUT: fake_bl_100 
* OUTPUT: fake_br_100 
* OUTPUT: fake_bl_101 
* OUTPUT: fake_br_101 
* OUTPUT: fake_bl_102 
* OUTPUT: fake_br_102 
* OUTPUT: fake_bl_103 
* OUTPUT: fake_br_103 
* OUTPUT: fake_bl_104 
* OUTPUT: fake_br_104 
* OUTPUT: fake_bl_105 
* OUTPUT: fake_br_105 
* OUTPUT: fake_bl_106 
* OUTPUT: fake_br_106 
* OUTPUT: fake_bl_107 
* OUTPUT: fake_br_107 
* OUTPUT: fake_bl_108 
* OUTPUT: fake_br_108 
* OUTPUT: fake_bl_109 
* OUTPUT: fake_br_109 
* OUTPUT: fake_bl_110 
* OUTPUT: fake_br_110 
* OUTPUT: fake_bl_111 
* OUTPUT: fake_br_111 
* OUTPUT: fake_bl_112 
* OUTPUT: fake_br_112 
* OUTPUT: fake_bl_113 
* OUTPUT: fake_br_113 
* OUTPUT: fake_bl_114 
* OUTPUT: fake_br_114 
* OUTPUT: fake_bl_115 
* OUTPUT: fake_br_115 
* OUTPUT: fake_bl_116 
* OUTPUT: fake_br_116 
* OUTPUT: fake_bl_117 
* OUTPUT: fake_br_117 
* OUTPUT: fake_bl_118 
* OUTPUT: fake_br_118 
* OUTPUT: fake_bl_119 
* OUTPUT: fake_br_119 
* OUTPUT: fake_bl_120 
* OUTPUT: fake_br_120 
* OUTPUT: fake_bl_121 
* OUTPUT: fake_br_121 
* OUTPUT: fake_bl_122 
* OUTPUT: fake_br_122 
* OUTPUT: fake_bl_123 
* OUTPUT: fake_br_123 
* OUTPUT: fake_bl_124 
* OUTPUT: fake_br_124 
* OUTPUT: fake_bl_125 
* OUTPUT: fake_br_125 
* OUTPUT: fake_bl_126 
* OUTPUT: fake_br_126 
* OUTPUT: fake_bl_127 
* OUTPUT: fake_br_127 
* OUTPUT: fake_bl_128 
* OUTPUT: fake_br_128 
* POWER : vdd 
* GROUND: gnd 
* BIAS  : gate 
Xrca_bottom_0
+ fake_bl_0 vdd gnd fake_br_0 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_1
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_2
+ fake_bl_1 vdd gnd fake_br_1 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_3
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_4
+ fake_bl_2 vdd gnd fake_br_2 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_5
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_6
+ fake_bl_3 vdd gnd fake_br_3 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_7
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_8
+ fake_bl_4 vdd gnd fake_br_4 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_9
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_10
+ fake_bl_5 vdd gnd fake_br_5 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_11
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_12
+ fake_bl_6 vdd gnd fake_br_6 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_13
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_14
+ fake_bl_7 vdd gnd fake_br_7 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_15
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_16
+ fake_bl_8 vdd gnd fake_br_8 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_17
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_18
+ fake_bl_9 vdd gnd fake_br_9 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_19
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_20
+ fake_bl_10 vdd gnd fake_br_10 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_21
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_22
+ fake_bl_11 vdd gnd fake_br_11 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_23
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_24
+ fake_bl_12 vdd gnd fake_br_12 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_25
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_26
+ fake_bl_13 vdd gnd fake_br_13 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_27
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_28
+ fake_bl_14 vdd gnd fake_br_14 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_29
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_30
+ fake_bl_15 vdd gnd fake_br_15 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_31
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_32
+ fake_bl_16 vdd gnd fake_br_16 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_33
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_34
+ fake_bl_17 vdd gnd fake_br_17 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_35
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_36
+ fake_bl_18 vdd gnd fake_br_18 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_37
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_38
+ fake_bl_19 vdd gnd fake_br_19 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_39
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_40
+ fake_bl_20 vdd gnd fake_br_20 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_41
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_42
+ fake_bl_21 vdd gnd fake_br_21 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_43
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_44
+ fake_bl_22 vdd gnd fake_br_22 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_45
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_46
+ fake_bl_23 vdd gnd fake_br_23 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_47
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_48
+ fake_bl_24 vdd gnd fake_br_24 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_49
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_50
+ fake_bl_25 vdd gnd fake_br_25 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_51
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_52
+ fake_bl_26 vdd gnd fake_br_26 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_53
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_54
+ fake_bl_27 vdd gnd fake_br_27 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_55
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_56
+ fake_bl_28 vdd gnd fake_br_28 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_57
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_58
+ fake_bl_29 vdd gnd fake_br_29 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_59
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_60
+ fake_bl_30 vdd gnd fake_br_30 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_61
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_62
+ fake_bl_31 vdd gnd fake_br_31 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_63
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_64
+ fake_bl_32 vdd gnd fake_br_32 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_65
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_66
+ fake_bl_33 vdd gnd fake_br_33 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_67
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_68
+ fake_bl_34 vdd gnd fake_br_34 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_69
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_70
+ fake_bl_35 vdd gnd fake_br_35 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_71
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_72
+ fake_bl_36 vdd gnd fake_br_36 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_73
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_74
+ fake_bl_37 vdd gnd fake_br_37 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_75
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_76
+ fake_bl_38 vdd gnd fake_br_38 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_77
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_78
+ fake_bl_39 vdd gnd fake_br_39 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_79
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_80
+ fake_bl_40 vdd gnd fake_br_40 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_81
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_82
+ fake_bl_41 vdd gnd fake_br_41 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_83
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_84
+ fake_bl_42 vdd gnd fake_br_42 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_85
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_86
+ fake_bl_43 vdd gnd fake_br_43 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_87
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_88
+ fake_bl_44 vdd gnd fake_br_44 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_89
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_90
+ fake_bl_45 vdd gnd fake_br_45 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_91
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_92
+ fake_bl_46 vdd gnd fake_br_46 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_93
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_94
+ fake_bl_47 vdd gnd fake_br_47 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_95
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_96
+ fake_bl_48 vdd gnd fake_br_48 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_97
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_98
+ fake_bl_49 vdd gnd fake_br_49 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_99
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_100
+ fake_bl_50 vdd gnd fake_br_50 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_101
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_102
+ fake_bl_51 vdd gnd fake_br_51 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_103
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_104
+ fake_bl_52 vdd gnd fake_br_52 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_105
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_106
+ fake_bl_53 vdd gnd fake_br_53 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_107
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_108
+ fake_bl_54 vdd gnd fake_br_54 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_109
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_110
+ fake_bl_55 vdd gnd fake_br_55 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_111
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_112
+ fake_bl_56 vdd gnd fake_br_56 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_113
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_114
+ fake_bl_57 vdd gnd fake_br_57 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_115
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_116
+ fake_bl_58 vdd gnd fake_br_58 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_117
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_118
+ fake_bl_59 vdd gnd fake_br_59 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_119
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_120
+ fake_bl_60 vdd gnd fake_br_60 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_121
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_122
+ fake_bl_61 vdd gnd fake_br_61 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_123
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_124
+ fake_bl_62 vdd gnd fake_br_62 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_125
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_126
+ fake_bl_63 vdd gnd fake_br_63 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_127
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_128
+ fake_bl_64 vdd gnd fake_br_64 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_129
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_130
+ fake_bl_65 vdd gnd fake_br_65 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_131
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_132
+ fake_bl_66 vdd gnd fake_br_66 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_133
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_134
+ fake_bl_67 vdd gnd fake_br_67 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_135
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_136
+ fake_bl_68 vdd gnd fake_br_68 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_137
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_138
+ fake_bl_69 vdd gnd fake_br_69 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_139
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_140
+ fake_bl_70 vdd gnd fake_br_70 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_141
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_142
+ fake_bl_71 vdd gnd fake_br_71 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_143
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_144
+ fake_bl_72 vdd gnd fake_br_72 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_145
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_146
+ fake_bl_73 vdd gnd fake_br_73 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_147
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_148
+ fake_bl_74 vdd gnd fake_br_74 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_149
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_150
+ fake_bl_75 vdd gnd fake_br_75 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_151
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_152
+ fake_bl_76 vdd gnd fake_br_76 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_153
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_154
+ fake_bl_77 vdd gnd fake_br_77 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_155
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_156
+ fake_bl_78 vdd gnd fake_br_78 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_157
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_158
+ fake_bl_79 vdd gnd fake_br_79 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_159
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_160
+ fake_bl_80 vdd gnd fake_br_80 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_161
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_162
+ fake_bl_81 vdd gnd fake_br_81 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_163
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_164
+ fake_bl_82 vdd gnd fake_br_82 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_165
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_166
+ fake_bl_83 vdd gnd fake_br_83 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_167
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_168
+ fake_bl_84 vdd gnd fake_br_84 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_169
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_170
+ fake_bl_85 vdd gnd fake_br_85 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_171
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_172
+ fake_bl_86 vdd gnd fake_br_86 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_173
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_174
+ fake_bl_87 vdd gnd fake_br_87 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_175
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_176
+ fake_bl_88 vdd gnd fake_br_88 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_177
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_178
+ fake_bl_89 vdd gnd fake_br_89 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_179
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_180
+ fake_bl_90 vdd gnd fake_br_90 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_181
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_182
+ fake_bl_91 vdd gnd fake_br_91 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_183
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_184
+ fake_bl_92 vdd gnd fake_br_92 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_185
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_186
+ fake_bl_93 vdd gnd fake_br_93 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_187
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_188
+ fake_bl_94 vdd gnd fake_br_94 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_189
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_190
+ fake_bl_95 vdd gnd fake_br_95 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_191
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_192
+ fake_bl_96 vdd gnd fake_br_96 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_193
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_194
+ fake_bl_97 vdd gnd fake_br_97 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_195
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_196
+ fake_bl_98 vdd gnd fake_br_98 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_197
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_198
+ fake_bl_99 vdd gnd fake_br_99 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_199
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_200
+ fake_bl_100 vdd gnd fake_br_100 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_201
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_202
+ fake_bl_101 vdd gnd fake_br_101 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_203
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_204
+ fake_bl_102 vdd gnd fake_br_102 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_205
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_206
+ fake_bl_103 vdd gnd fake_br_103 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_207
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_208
+ fake_bl_104 vdd gnd fake_br_104 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_209
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_210
+ fake_bl_105 vdd gnd fake_br_105 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_211
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_212
+ fake_bl_106 vdd gnd fake_br_106 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_213
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_214
+ fake_bl_107 vdd gnd fake_br_107 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_215
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_216
+ fake_bl_108 vdd gnd fake_br_108 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_217
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_218
+ fake_bl_109 vdd gnd fake_br_109 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_219
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_220
+ fake_bl_110 vdd gnd fake_br_110 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_221
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_222
+ fake_bl_111 vdd gnd fake_br_111 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_223
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_224
+ fake_bl_112 vdd gnd fake_br_112 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_225
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_226
+ fake_bl_113 vdd gnd fake_br_113 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_227
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_228
+ fake_bl_114 vdd gnd fake_br_114 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_229
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_230
+ fake_bl_115 vdd gnd fake_br_115 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_231
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_232
+ fake_bl_116 vdd gnd fake_br_116 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_233
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_234
+ fake_bl_117 vdd gnd fake_br_117 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_235
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_236
+ fake_bl_118 vdd gnd fake_br_118 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_237
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_238
+ fake_bl_119 vdd gnd fake_br_119 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_239
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_240
+ fake_bl_120 vdd gnd fake_br_120 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_241
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_242
+ fake_bl_121 vdd gnd fake_br_121 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_243
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_244
+ fake_bl_122 vdd gnd fake_br_122 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_245
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_246
+ fake_bl_123 vdd gnd fake_br_123 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_247
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_248
+ fake_bl_124 vdd gnd fake_br_124 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_249
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_250
+ fake_bl_125 vdd gnd fake_br_125 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_251
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_252
+ fake_bl_126 vdd gnd fake_br_126 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_253
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda_cent
Xrca_bottom_254
+ fake_bl_127 vdd gnd fake_br_127 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
Xrca_bottom_255
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colenda_p_cent
Xrca_bottom_256
+ fake_bl_128 vdd gnd fake_br_128 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colenda
.ENDS sky130_sram_1kbyte_1rw_32x256_8_sky130_col_cap_array_0
* NGSPICE file created from sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy BL BR VGND VPWR VPB VNB WL
X0 ll WL BR VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
X1 ul Q_bar_float VGND VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
X2 BL WL ul VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
*X3 ur WL ur VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
*X4 lr WL lr VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
X5 VPWR Q_float lr VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X6 ur Q_bar_float VPWR VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X7 VGND Q_float ll VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_wlstrapa.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_wlstrapa VPWR
.ends

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_sky130_dummy_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 wl_0_0 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INPUT : wl_0_0 
* POWER : vdd 
* GROUND: gnd 
Xrow_0_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_0_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
Xrow_0_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_0_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__openram_sp_cell_opt1a_dummy
.ENDS sky130_sram_1kbyte_1rw_32x256_8_sky130_dummy_array
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_rowend.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_rowend VPWR WL
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_rowenda.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_rowenda VPWR WL
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_cornerb.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_cornerb VPWR VPB VNB
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_cornera.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_cornera VNB VPWR VPB
.ends

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_sky130_row_cap_array_0
+ wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9
+ wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17
+ wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25
+ wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33
+ wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41
+ wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49
+ wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57
+ wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65
+ wl_0_66 wl_0_67 vdd gnd
* OUTPUT: wl_0_0 
* OUTPUT: wl_0_1 
* OUTPUT: wl_0_2 
* OUTPUT: wl_0_3 
* OUTPUT: wl_0_4 
* OUTPUT: wl_0_5 
* OUTPUT: wl_0_6 
* OUTPUT: wl_0_7 
* OUTPUT: wl_0_8 
* OUTPUT: wl_0_9 
* OUTPUT: wl_0_10 
* OUTPUT: wl_0_11 
* OUTPUT: wl_0_12 
* OUTPUT: wl_0_13 
* OUTPUT: wl_0_14 
* OUTPUT: wl_0_15 
* OUTPUT: wl_0_16 
* OUTPUT: wl_0_17 
* OUTPUT: wl_0_18 
* OUTPUT: wl_0_19 
* OUTPUT: wl_0_20 
* OUTPUT: wl_0_21 
* OUTPUT: wl_0_22 
* OUTPUT: wl_0_23 
* OUTPUT: wl_0_24 
* OUTPUT: wl_0_25 
* OUTPUT: wl_0_26 
* OUTPUT: wl_0_27 
* OUTPUT: wl_0_28 
* OUTPUT: wl_0_29 
* OUTPUT: wl_0_30 
* OUTPUT: wl_0_31 
* OUTPUT: wl_0_32 
* OUTPUT: wl_0_33 
* OUTPUT: wl_0_34 
* OUTPUT: wl_0_35 
* OUTPUT: wl_0_36 
* OUTPUT: wl_0_37 
* OUTPUT: wl_0_38 
* OUTPUT: wl_0_39 
* OUTPUT: wl_0_40 
* OUTPUT: wl_0_41 
* OUTPUT: wl_0_42 
* OUTPUT: wl_0_43 
* OUTPUT: wl_0_44 
* OUTPUT: wl_0_45 
* OUTPUT: wl_0_46 
* OUTPUT: wl_0_47 
* OUTPUT: wl_0_48 
* OUTPUT: wl_0_49 
* OUTPUT: wl_0_50 
* OUTPUT: wl_0_51 
* OUTPUT: wl_0_52 
* OUTPUT: wl_0_53 
* OUTPUT: wl_0_54 
* OUTPUT: wl_0_55 
* OUTPUT: wl_0_56 
* OUTPUT: wl_0_57 
* OUTPUT: wl_0_58 
* OUTPUT: wl_0_59 
* OUTPUT: wl_0_60 
* OUTPUT: wl_0_61 
* OUTPUT: wl_0_62 
* OUTPUT: wl_0_63 
* OUTPUT: wl_0_64 
* OUTPUT: wl_0_65 
* OUTPUT: wl_0_66 
* OUTPUT: wl_0_67 
* POWER : vdd 
* GROUND: gnd 
Xrca_0
+ vdd gnd vdd
+ sky130_fd_bd_sram__sram_sp_cornera
Xrca_1
+ wl_0_0 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_2
+ wl_0_1 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_3
+ wl_0_2 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_4
+ wl_0_3 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_5
+ wl_0_4 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_6
+ wl_0_5 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_7
+ wl_0_6 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_8
+ wl_0_7 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_9
+ wl_0_8 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_10
+ wl_0_9 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_11
+ wl_0_10 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_12
+ wl_0_11 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_13
+ wl_0_12 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_14
+ wl_0_13 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_15
+ wl_0_14 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_16
+ wl_0_15 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_17
+ wl_0_16 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_18
+ wl_0_17 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_19
+ wl_0_18 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_20
+ wl_0_19 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_21
+ wl_0_20 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_22
+ wl_0_21 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_23
+ wl_0_22 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_24
+ wl_0_23 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_25
+ wl_0_24 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_26
+ wl_0_25 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_27
+ wl_0_26 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_28
+ wl_0_27 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_29
+ wl_0_28 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_30
+ wl_0_29 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_31
+ wl_0_30 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_32
+ wl_0_31 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_33
+ wl_0_32 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_34
+ wl_0_33 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_35
+ wl_0_34 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_36
+ wl_0_35 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_37
+ wl_0_36 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_38
+ wl_0_37 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_39
+ wl_0_38 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_40
+ wl_0_39 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_41
+ wl_0_40 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_42
+ wl_0_41 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_43
+ wl_0_42 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_44
+ wl_0_43 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_45
+ wl_0_44 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_46
+ wl_0_45 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_47
+ wl_0_46 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_48
+ wl_0_47 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_49
+ wl_0_48 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_50
+ wl_0_49 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_51
+ wl_0_50 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_52
+ wl_0_51 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_53
+ wl_0_52 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_54
+ wl_0_53 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_55
+ wl_0_54 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_56
+ wl_0_55 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_57
+ wl_0_56 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_58
+ wl_0_57 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_59
+ wl_0_58 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_60
+ wl_0_59 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_61
+ wl_0_60 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_62
+ wl_0_61 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_63
+ wl_0_62 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_64
+ wl_0_63 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_65
+ wl_0_64 vdd
+ sky130_fd_bd_sram__sram_sp_rowenda
Xrca_66
+ wl_0_65 vdd
+ sky130_fd_bd_sram__sram_sp_rowend
Xrca_67
+ vdd gnd vdd
+ sky130_fd_bd_sram__sram_sp_cornerb
.ENDS sky130_sram_1kbyte_1rw_32x256_8_sky130_row_cap_array_0
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_cell_opt1a.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_cell_opt1a BL BR VGND VPWR VPB VNB WL
X0 Q_bar WL BR VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
X1 Q Q_bar VGND VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
*X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
*X4 Q_bar WL Q_bar VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
X5 VPWR Q Q_bar VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X6 Q Q_bar VPWR VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X7 VGND Q Q_bar VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_cell_opt1.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_cell_opt1 BL BR VGND VPWR VPB VNB WL
X0 Q_bar WL BR VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
X1 Q Q_bar VGND VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass w=0.14 l=0.15
*X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
*X4 Q_bar WL Q_bar VPB sky130_fd_pr__special_pfet_pass w=0.07 l=0.095
X5 VPWR Q Q_bar VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X6 Q Q_bar VPWR VPB sky130_fd_pr__special_pfet_pass w=0.14 l=0.15
X7 VGND Q Q_bar VNB sky130_fd_pr__special_nfet_latch w=0.21 l=0.15
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_wlstrap.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_wlstrap VPWR
.ends

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_sky130_bitcell_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 wl_0_0 wl_0_1 wl_0_2
+ wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11
+ wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19
+ wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27
+ wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35
+ wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43
+ wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51
+ wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59
+ wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* POWER : vdd 
* GROUND: gnd 
* rows: 65 cols: 129
Xrow_0_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_0_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_0_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_0_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_0
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_1_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_1_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_1_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_1_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_1
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_2_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_2_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_2_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_2_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_2
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_3_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_3_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_3_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_3_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_3
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_4_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_4_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_4_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_4_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_4
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_5_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_5_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_5_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_5_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_5
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_6_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_6_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_6_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_6_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_6
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_7_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_7_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_7_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_7_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_7
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_8_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_8_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_8_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_8_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_8
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_9_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_9_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_9_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_9_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_9
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_10_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_10_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_10_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_10_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_10
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_11_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_11_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_11_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_11_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_11
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_12_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_12_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_12_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_12_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_12
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_13_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_13_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_13_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_13_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_13
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_14_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_14_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_14_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_14_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_14
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_15_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_15_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_15_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_15_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_15
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_16_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_16_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_16_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_16_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_16
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_17_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_17_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_17_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_17_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_17
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_18_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_18_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_18_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_18_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_18
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_19_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_19_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_19_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_19_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_19
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_20_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_20_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_20_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_20_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_20
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_21_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_21_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_21_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_21_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_21
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_22_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_22_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_22_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_22_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_22
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_23_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_23_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_23_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_23_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_23
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_24_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_24_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_24_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_24_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_24
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_25_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_25_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_25_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_25_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_25
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_26_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_26_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_26_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_26_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_26
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_27_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_27_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_27_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_27_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_27
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_28_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_28_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_28_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_28_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_28
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_29_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_29_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_29_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_29_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_29
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_30_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_30_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_30_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_30_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_30
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_31_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_31_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_31_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_31_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_31
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_32_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_32_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_32_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_32_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_32
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_33_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_33_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_33_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_33_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_33
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_34_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_34_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_34_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_34_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_34
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_35_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_35_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_35_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_35_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_35
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_36_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_36_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_36_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_36_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_36
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_37_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_37_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_37_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_37_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_37
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_38_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_38_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_38_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_38_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_38
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_39_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_39_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_39_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_39_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_39
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_40_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_40_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_40_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_40_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_40
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_41_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_41_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_41_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_41_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_41
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_42_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_42_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_42_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_42_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_42
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_43_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_43_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_43_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_43_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_43
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_44_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_44_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_44_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_44_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_44
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_45_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_45_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_45_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_45_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_45
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_46_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_46_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_46_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_46_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_46
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_47_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_47_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_47_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_47_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_47
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_48_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_48_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_48_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_48_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_48
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_49_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_49_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_49_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_49_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_49
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_50_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_50_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_50_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_50_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_50
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_51_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_51_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_51_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_51_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_51
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_52_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_52_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_52_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_52_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_52
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_53_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_53_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_53_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_53_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_53
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_54_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_54_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_54_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_54_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_54
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_55_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_55_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_55_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_55_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_55
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_56_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_56_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_56_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_56_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_56
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_57_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_57_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_57_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_57_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_57
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_58_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_58_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_58_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_58_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_58
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_59_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_59_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_59_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_59_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_59
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_60_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_60_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_60_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_60_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_60
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_61_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_61_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_61_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_61_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_61
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_62_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_62_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_62_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_62_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_62
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_63_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_0_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_1_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_2_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_3_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_4_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_5_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_6_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_7_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_8_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_9_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_10_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_11_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_12_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_13_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_14_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_15_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_16_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_17_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_18_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_19_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_20_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_21_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_22_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_23_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_24_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_25_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_26_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_27_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_28_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_29_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_30_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_31_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_32_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_33_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_34_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_35_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_36_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_37_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_38_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_39_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_40_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_41_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_42_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_43_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_44_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_45_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_46_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_47_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_48_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_49_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_50_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_51_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_52_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_53_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_54_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_55_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_56_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_57_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_58_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_59_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_60_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_61_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_62_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_63_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_64_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_65_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_66_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_67_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_68_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_69_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_70_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_71_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_72_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_73_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_74_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_75_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_76_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_77_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_78_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_79_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_80_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_81_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_82_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_83_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_84_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_85_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_86_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_87_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_88_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_89_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_90_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_91_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_92_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_93_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_94_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_95_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_96_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_97_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_98_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_99_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_100_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_101_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_102_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_103_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_104_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_105_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_106_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_107_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_108_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_109_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_110_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_111_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_112_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_113_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_114_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_115_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_116_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_117_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_118_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_119_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_120_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_121_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_122_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_123_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_124_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_125_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_126_wlstrapa
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrapa
Xrow_63_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_63_col_127_wlstrapa_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrapa_p
Xrow_63_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_63
+ sky130_fd_bd_sram__sram_sp_cell_opt1a
Xrow_64_col_0_bitcell
+ bl_0_0 br_0_0 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_0_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_1_bitcell
+ bl_0_1 br_0_1 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_1_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_2_bitcell
+ bl_0_2 br_0_2 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_2_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_3_bitcell
+ bl_0_3 br_0_3 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_3_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_4_bitcell
+ bl_0_4 br_0_4 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_4_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_5_bitcell
+ bl_0_5 br_0_5 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_5_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_6_bitcell
+ bl_0_6 br_0_6 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_6_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_7_bitcell
+ bl_0_7 br_0_7 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_7_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_8_bitcell
+ bl_0_8 br_0_8 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_8_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_9_bitcell
+ bl_0_9 br_0_9 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_9_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_10_bitcell
+ bl_0_10 br_0_10 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_10_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_11_bitcell
+ bl_0_11 br_0_11 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_11_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_12_bitcell
+ bl_0_12 br_0_12 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_12_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_13_bitcell
+ bl_0_13 br_0_13 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_13_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_14_bitcell
+ bl_0_14 br_0_14 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_14_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_15_bitcell
+ bl_0_15 br_0_15 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_15_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_16_bitcell
+ bl_0_16 br_0_16 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_16_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_17_bitcell
+ bl_0_17 br_0_17 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_17_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_18_bitcell
+ bl_0_18 br_0_18 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_18_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_19_bitcell
+ bl_0_19 br_0_19 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_19_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_20_bitcell
+ bl_0_20 br_0_20 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_20_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_21_bitcell
+ bl_0_21 br_0_21 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_21_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_22_bitcell
+ bl_0_22 br_0_22 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_22_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_23_bitcell
+ bl_0_23 br_0_23 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_23_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_24_bitcell
+ bl_0_24 br_0_24 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_24_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_25_bitcell
+ bl_0_25 br_0_25 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_25_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_26_bitcell
+ bl_0_26 br_0_26 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_26_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_27_bitcell
+ bl_0_27 br_0_27 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_27_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_28_bitcell
+ bl_0_28 br_0_28 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_28_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_29_bitcell
+ bl_0_29 br_0_29 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_29_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_30_bitcell
+ bl_0_30 br_0_30 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_30_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_31_bitcell
+ bl_0_31 br_0_31 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_31_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_32_bitcell
+ bl_0_32 br_0_32 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_32_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_33_bitcell
+ bl_0_33 br_0_33 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_33_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_34_bitcell
+ bl_0_34 br_0_34 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_34_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_35_bitcell
+ bl_0_35 br_0_35 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_35_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_36_bitcell
+ bl_0_36 br_0_36 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_36_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_37_bitcell
+ bl_0_37 br_0_37 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_37_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_38_bitcell
+ bl_0_38 br_0_38 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_38_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_39_bitcell
+ bl_0_39 br_0_39 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_39_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_40_bitcell
+ bl_0_40 br_0_40 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_40_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_41_bitcell
+ bl_0_41 br_0_41 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_41_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_42_bitcell
+ bl_0_42 br_0_42 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_42_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_43_bitcell
+ bl_0_43 br_0_43 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_43_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_44_bitcell
+ bl_0_44 br_0_44 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_44_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_45_bitcell
+ bl_0_45 br_0_45 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_45_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_46_bitcell
+ bl_0_46 br_0_46 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_46_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_47_bitcell
+ bl_0_47 br_0_47 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_47_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_48_bitcell
+ bl_0_48 br_0_48 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_48_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_49_bitcell
+ bl_0_49 br_0_49 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_49_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_50_bitcell
+ bl_0_50 br_0_50 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_50_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_51_bitcell
+ bl_0_51 br_0_51 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_51_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_52_bitcell
+ bl_0_52 br_0_52 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_52_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_53_bitcell
+ bl_0_53 br_0_53 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_53_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_54_bitcell
+ bl_0_54 br_0_54 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_54_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_55_bitcell
+ bl_0_55 br_0_55 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_55_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_56_bitcell
+ bl_0_56 br_0_56 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_56_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_57_bitcell
+ bl_0_57 br_0_57 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_57_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_58_bitcell
+ bl_0_58 br_0_58 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_58_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_59_bitcell
+ bl_0_59 br_0_59 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_59_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_60_bitcell
+ bl_0_60 br_0_60 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_60_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_61_bitcell
+ bl_0_61 br_0_61 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_61_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_62_bitcell
+ bl_0_62 br_0_62 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_62_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_63_bitcell
+ bl_0_63 br_0_63 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_63_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_64_bitcell
+ bl_0_64 br_0_64 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_64_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_65_bitcell
+ bl_0_65 br_0_65 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_65_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_66_bitcell
+ bl_0_66 br_0_66 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_66_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_67_bitcell
+ bl_0_67 br_0_67 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_67_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_68_bitcell
+ bl_0_68 br_0_68 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_68_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_69_bitcell
+ bl_0_69 br_0_69 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_69_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_70_bitcell
+ bl_0_70 br_0_70 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_70_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_71_bitcell
+ bl_0_71 br_0_71 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_71_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_72_bitcell
+ bl_0_72 br_0_72 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_72_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_73_bitcell
+ bl_0_73 br_0_73 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_73_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_74_bitcell
+ bl_0_74 br_0_74 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_74_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_75_bitcell
+ bl_0_75 br_0_75 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_75_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_76_bitcell
+ bl_0_76 br_0_76 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_76_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_77_bitcell
+ bl_0_77 br_0_77 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_77_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_78_bitcell
+ bl_0_78 br_0_78 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_78_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_79_bitcell
+ bl_0_79 br_0_79 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_79_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_80_bitcell
+ bl_0_80 br_0_80 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_80_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_81_bitcell
+ bl_0_81 br_0_81 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_81_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_82_bitcell
+ bl_0_82 br_0_82 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_82_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_83_bitcell
+ bl_0_83 br_0_83 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_83_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_84_bitcell
+ bl_0_84 br_0_84 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_84_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_85_bitcell
+ bl_0_85 br_0_85 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_85_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_86_bitcell
+ bl_0_86 br_0_86 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_86_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_87_bitcell
+ bl_0_87 br_0_87 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_87_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_88_bitcell
+ bl_0_88 br_0_88 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_88_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_89_bitcell
+ bl_0_89 br_0_89 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_89_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_90_bitcell
+ bl_0_90 br_0_90 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_90_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_91_bitcell
+ bl_0_91 br_0_91 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_91_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_92_bitcell
+ bl_0_92 br_0_92 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_92_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_93_bitcell
+ bl_0_93 br_0_93 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_93_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_94_bitcell
+ bl_0_94 br_0_94 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_94_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_95_bitcell
+ bl_0_95 br_0_95 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_95_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_96_bitcell
+ bl_0_96 br_0_96 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_96_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_97_bitcell
+ bl_0_97 br_0_97 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_97_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_98_bitcell
+ bl_0_98 br_0_98 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_98_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_99_bitcell
+ bl_0_99 br_0_99 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_99_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_100_bitcell
+ bl_0_100 br_0_100 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_100_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_101_bitcell
+ bl_0_101 br_0_101 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_101_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_102_bitcell
+ bl_0_102 br_0_102 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_102_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_103_bitcell
+ bl_0_103 br_0_103 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_103_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_104_bitcell
+ bl_0_104 br_0_104 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_104_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_105_bitcell
+ bl_0_105 br_0_105 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_105_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_106_bitcell
+ bl_0_106 br_0_106 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_106_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_107_bitcell
+ bl_0_107 br_0_107 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_107_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_108_bitcell
+ bl_0_108 br_0_108 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_108_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_109_bitcell
+ bl_0_109 br_0_109 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_109_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_110_bitcell
+ bl_0_110 br_0_110 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_110_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_111_bitcell
+ bl_0_111 br_0_111 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_111_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_112_bitcell
+ bl_0_112 br_0_112 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_112_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_113_bitcell
+ bl_0_113 br_0_113 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_113_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_114_bitcell
+ bl_0_114 br_0_114 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_114_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_115_bitcell
+ bl_0_115 br_0_115 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_115_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_116_bitcell
+ bl_0_116 br_0_116 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_116_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_117_bitcell
+ bl_0_117 br_0_117 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_117_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_118_bitcell
+ bl_0_118 br_0_118 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_118_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_119_bitcell
+ bl_0_119 br_0_119 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_119_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_120_bitcell
+ bl_0_120 br_0_120 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_120_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_121_bitcell
+ bl_0_121 br_0_121 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_121_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_122_bitcell
+ bl_0_122 br_0_122 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_122_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_123_bitcell
+ bl_0_123 br_0_123 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_123_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_124_bitcell
+ bl_0_124 br_0_124 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_124_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_125_bitcell
+ bl_0_125 br_0_125 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_125_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_126_bitcell
+ bl_0_126 br_0_126 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_126_wlstrap
+ vdd
+ sky130_fd_bd_sram__sram_sp_wlstrap
Xrow_64_col_127_bitcell
+ bl_0_127 br_0_127 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
Xrow_64_col_127_wlstrap_p
+ gnd
+ sky130_fd_bd_sram__sram_sp_wlstrap_p
Xrow_64_col_128_bitcell
+ bl_0_128 br_0_128 gnd vdd vdd gnd wl_0_64
+ sky130_fd_bd_sram__sram_sp_cell_opt1
.ENDS sky130_sram_1kbyte_1rw_32x256_8_sky130_bitcell_array
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_colend_cent.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_colend_cent VPWR VPB VNB
.ends

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_sky130_col_cap_array
+ fake_bl_0 fake_br_0 fake_bl_1 fake_br_1 fake_bl_2 fake_br_2 fake_bl_3
+ fake_br_3 fake_bl_4 fake_br_4 fake_bl_5 fake_br_5 fake_bl_6 fake_br_6
+ fake_bl_7 fake_br_7 fake_bl_8 fake_br_8 fake_bl_9 fake_br_9 fake_bl_10
+ fake_br_10 fake_bl_11 fake_br_11 fake_bl_12 fake_br_12 fake_bl_13
+ fake_br_13 fake_bl_14 fake_br_14 fake_bl_15 fake_br_15 fake_bl_16
+ fake_br_16 fake_bl_17 fake_br_17 fake_bl_18 fake_br_18 fake_bl_19
+ fake_br_19 fake_bl_20 fake_br_20 fake_bl_21 fake_br_21 fake_bl_22
+ fake_br_22 fake_bl_23 fake_br_23 fake_bl_24 fake_br_24 fake_bl_25
+ fake_br_25 fake_bl_26 fake_br_26 fake_bl_27 fake_br_27 fake_bl_28
+ fake_br_28 fake_bl_29 fake_br_29 fake_bl_30 fake_br_30 fake_bl_31
+ fake_br_31 fake_bl_32 fake_br_32 fake_bl_33 fake_br_33 fake_bl_34
+ fake_br_34 fake_bl_35 fake_br_35 fake_bl_36 fake_br_36 fake_bl_37
+ fake_br_37 fake_bl_38 fake_br_38 fake_bl_39 fake_br_39 fake_bl_40
+ fake_br_40 fake_bl_41 fake_br_41 fake_bl_42 fake_br_42 fake_bl_43
+ fake_br_43 fake_bl_44 fake_br_44 fake_bl_45 fake_br_45 fake_bl_46
+ fake_br_46 fake_bl_47 fake_br_47 fake_bl_48 fake_br_48 fake_bl_49
+ fake_br_49 fake_bl_50 fake_br_50 fake_bl_51 fake_br_51 fake_bl_52
+ fake_br_52 fake_bl_53 fake_br_53 fake_bl_54 fake_br_54 fake_bl_55
+ fake_br_55 fake_bl_56 fake_br_56 fake_bl_57 fake_br_57 fake_bl_58
+ fake_br_58 fake_bl_59 fake_br_59 fake_bl_60 fake_br_60 fake_bl_61
+ fake_br_61 fake_bl_62 fake_br_62 fake_bl_63 fake_br_63 fake_bl_64
+ fake_br_64 fake_bl_65 fake_br_65 fake_bl_66 fake_br_66 fake_bl_67
+ fake_br_67 fake_bl_68 fake_br_68 fake_bl_69 fake_br_69 fake_bl_70
+ fake_br_70 fake_bl_71 fake_br_71 fake_bl_72 fake_br_72 fake_bl_73
+ fake_br_73 fake_bl_74 fake_br_74 fake_bl_75 fake_br_75 fake_bl_76
+ fake_br_76 fake_bl_77 fake_br_77 fake_bl_78 fake_br_78 fake_bl_79
+ fake_br_79 fake_bl_80 fake_br_80 fake_bl_81 fake_br_81 fake_bl_82
+ fake_br_82 fake_bl_83 fake_br_83 fake_bl_84 fake_br_84 fake_bl_85
+ fake_br_85 fake_bl_86 fake_br_86 fake_bl_87 fake_br_87 fake_bl_88
+ fake_br_88 fake_bl_89 fake_br_89 fake_bl_90 fake_br_90 fake_bl_91
+ fake_br_91 fake_bl_92 fake_br_92 fake_bl_93 fake_br_93 fake_bl_94
+ fake_br_94 fake_bl_95 fake_br_95 fake_bl_96 fake_br_96 fake_bl_97
+ fake_br_97 fake_bl_98 fake_br_98 fake_bl_99 fake_br_99 fake_bl_100
+ fake_br_100 fake_bl_101 fake_br_101 fake_bl_102 fake_br_102
+ fake_bl_103 fake_br_103 fake_bl_104 fake_br_104 fake_bl_105
+ fake_br_105 fake_bl_106 fake_br_106 fake_bl_107 fake_br_107
+ fake_bl_108 fake_br_108 fake_bl_109 fake_br_109 fake_bl_110
+ fake_br_110 fake_bl_111 fake_br_111 fake_bl_112 fake_br_112
+ fake_bl_113 fake_br_113 fake_bl_114 fake_br_114 fake_bl_115
+ fake_br_115 fake_bl_116 fake_br_116 fake_bl_117 fake_br_117
+ fake_bl_118 fake_br_118 fake_bl_119 fake_br_119 fake_bl_120
+ fake_br_120 fake_bl_121 fake_br_121 fake_bl_122 fake_br_122
+ fake_bl_123 fake_br_123 fake_bl_124 fake_br_124 fake_bl_125
+ fake_br_125 fake_bl_126 fake_br_126 fake_bl_127 fake_br_127
+ fake_bl_128 fake_br_128 vdd gnd gate
* OUTPUT: fake_bl_0 
* OUTPUT: fake_br_0 
* OUTPUT: fake_bl_1 
* OUTPUT: fake_br_1 
* OUTPUT: fake_bl_2 
* OUTPUT: fake_br_2 
* OUTPUT: fake_bl_3 
* OUTPUT: fake_br_3 
* OUTPUT: fake_bl_4 
* OUTPUT: fake_br_4 
* OUTPUT: fake_bl_5 
* OUTPUT: fake_br_5 
* OUTPUT: fake_bl_6 
* OUTPUT: fake_br_6 
* OUTPUT: fake_bl_7 
* OUTPUT: fake_br_7 
* OUTPUT: fake_bl_8 
* OUTPUT: fake_br_8 
* OUTPUT: fake_bl_9 
* OUTPUT: fake_br_9 
* OUTPUT: fake_bl_10 
* OUTPUT: fake_br_10 
* OUTPUT: fake_bl_11 
* OUTPUT: fake_br_11 
* OUTPUT: fake_bl_12 
* OUTPUT: fake_br_12 
* OUTPUT: fake_bl_13 
* OUTPUT: fake_br_13 
* OUTPUT: fake_bl_14 
* OUTPUT: fake_br_14 
* OUTPUT: fake_bl_15 
* OUTPUT: fake_br_15 
* OUTPUT: fake_bl_16 
* OUTPUT: fake_br_16 
* OUTPUT: fake_bl_17 
* OUTPUT: fake_br_17 
* OUTPUT: fake_bl_18 
* OUTPUT: fake_br_18 
* OUTPUT: fake_bl_19 
* OUTPUT: fake_br_19 
* OUTPUT: fake_bl_20 
* OUTPUT: fake_br_20 
* OUTPUT: fake_bl_21 
* OUTPUT: fake_br_21 
* OUTPUT: fake_bl_22 
* OUTPUT: fake_br_22 
* OUTPUT: fake_bl_23 
* OUTPUT: fake_br_23 
* OUTPUT: fake_bl_24 
* OUTPUT: fake_br_24 
* OUTPUT: fake_bl_25 
* OUTPUT: fake_br_25 
* OUTPUT: fake_bl_26 
* OUTPUT: fake_br_26 
* OUTPUT: fake_bl_27 
* OUTPUT: fake_br_27 
* OUTPUT: fake_bl_28 
* OUTPUT: fake_br_28 
* OUTPUT: fake_bl_29 
* OUTPUT: fake_br_29 
* OUTPUT: fake_bl_30 
* OUTPUT: fake_br_30 
* OUTPUT: fake_bl_31 
* OUTPUT: fake_br_31 
* OUTPUT: fake_bl_32 
* OUTPUT: fake_br_32 
* OUTPUT: fake_bl_33 
* OUTPUT: fake_br_33 
* OUTPUT: fake_bl_34 
* OUTPUT: fake_br_34 
* OUTPUT: fake_bl_35 
* OUTPUT: fake_br_35 
* OUTPUT: fake_bl_36 
* OUTPUT: fake_br_36 
* OUTPUT: fake_bl_37 
* OUTPUT: fake_br_37 
* OUTPUT: fake_bl_38 
* OUTPUT: fake_br_38 
* OUTPUT: fake_bl_39 
* OUTPUT: fake_br_39 
* OUTPUT: fake_bl_40 
* OUTPUT: fake_br_40 
* OUTPUT: fake_bl_41 
* OUTPUT: fake_br_41 
* OUTPUT: fake_bl_42 
* OUTPUT: fake_br_42 
* OUTPUT: fake_bl_43 
* OUTPUT: fake_br_43 
* OUTPUT: fake_bl_44 
* OUTPUT: fake_br_44 
* OUTPUT: fake_bl_45 
* OUTPUT: fake_br_45 
* OUTPUT: fake_bl_46 
* OUTPUT: fake_br_46 
* OUTPUT: fake_bl_47 
* OUTPUT: fake_br_47 
* OUTPUT: fake_bl_48 
* OUTPUT: fake_br_48 
* OUTPUT: fake_bl_49 
* OUTPUT: fake_br_49 
* OUTPUT: fake_bl_50 
* OUTPUT: fake_br_50 
* OUTPUT: fake_bl_51 
* OUTPUT: fake_br_51 
* OUTPUT: fake_bl_52 
* OUTPUT: fake_br_52 
* OUTPUT: fake_bl_53 
* OUTPUT: fake_br_53 
* OUTPUT: fake_bl_54 
* OUTPUT: fake_br_54 
* OUTPUT: fake_bl_55 
* OUTPUT: fake_br_55 
* OUTPUT: fake_bl_56 
* OUTPUT: fake_br_56 
* OUTPUT: fake_bl_57 
* OUTPUT: fake_br_57 
* OUTPUT: fake_bl_58 
* OUTPUT: fake_br_58 
* OUTPUT: fake_bl_59 
* OUTPUT: fake_br_59 
* OUTPUT: fake_bl_60 
* OUTPUT: fake_br_60 
* OUTPUT: fake_bl_61 
* OUTPUT: fake_br_61 
* OUTPUT: fake_bl_62 
* OUTPUT: fake_br_62 
* OUTPUT: fake_bl_63 
* OUTPUT: fake_br_63 
* OUTPUT: fake_bl_64 
* OUTPUT: fake_br_64 
* OUTPUT: fake_bl_65 
* OUTPUT: fake_br_65 
* OUTPUT: fake_bl_66 
* OUTPUT: fake_br_66 
* OUTPUT: fake_bl_67 
* OUTPUT: fake_br_67 
* OUTPUT: fake_bl_68 
* OUTPUT: fake_br_68 
* OUTPUT: fake_bl_69 
* OUTPUT: fake_br_69 
* OUTPUT: fake_bl_70 
* OUTPUT: fake_br_70 
* OUTPUT: fake_bl_71 
* OUTPUT: fake_br_71 
* OUTPUT: fake_bl_72 
* OUTPUT: fake_br_72 
* OUTPUT: fake_bl_73 
* OUTPUT: fake_br_73 
* OUTPUT: fake_bl_74 
* OUTPUT: fake_br_74 
* OUTPUT: fake_bl_75 
* OUTPUT: fake_br_75 
* OUTPUT: fake_bl_76 
* OUTPUT: fake_br_76 
* OUTPUT: fake_bl_77 
* OUTPUT: fake_br_77 
* OUTPUT: fake_bl_78 
* OUTPUT: fake_br_78 
* OUTPUT: fake_bl_79 
* OUTPUT: fake_br_79 
* OUTPUT: fake_bl_80 
* OUTPUT: fake_br_80 
* OUTPUT: fake_bl_81 
* OUTPUT: fake_br_81 
* OUTPUT: fake_bl_82 
* OUTPUT: fake_br_82 
* OUTPUT: fake_bl_83 
* OUTPUT: fake_br_83 
* OUTPUT: fake_bl_84 
* OUTPUT: fake_br_84 
* OUTPUT: fake_bl_85 
* OUTPUT: fake_br_85 
* OUTPUT: fake_bl_86 
* OUTPUT: fake_br_86 
* OUTPUT: fake_bl_87 
* OUTPUT: fake_br_87 
* OUTPUT: fake_bl_88 
* OUTPUT: fake_br_88 
* OUTPUT: fake_bl_89 
* OUTPUT: fake_br_89 
* OUTPUT: fake_bl_90 
* OUTPUT: fake_br_90 
* OUTPUT: fake_bl_91 
* OUTPUT: fake_br_91 
* OUTPUT: fake_bl_92 
* OUTPUT: fake_br_92 
* OUTPUT: fake_bl_93 
* OUTPUT: fake_br_93 
* OUTPUT: fake_bl_94 
* OUTPUT: fake_br_94 
* OUTPUT: fake_bl_95 
* OUTPUT: fake_br_95 
* OUTPUT: fake_bl_96 
* OUTPUT: fake_br_96 
* OUTPUT: fake_bl_97 
* OUTPUT: fake_br_97 
* OUTPUT: fake_bl_98 
* OUTPUT: fake_br_98 
* OUTPUT: fake_bl_99 
* OUTPUT: fake_br_99 
* OUTPUT: fake_bl_100 
* OUTPUT: fake_br_100 
* OUTPUT: fake_bl_101 
* OUTPUT: fake_br_101 
* OUTPUT: fake_bl_102 
* OUTPUT: fake_br_102 
* OUTPUT: fake_bl_103 
* OUTPUT: fake_br_103 
* OUTPUT: fake_bl_104 
* OUTPUT: fake_br_104 
* OUTPUT: fake_bl_105 
* OUTPUT: fake_br_105 
* OUTPUT: fake_bl_106 
* OUTPUT: fake_br_106 
* OUTPUT: fake_bl_107 
* OUTPUT: fake_br_107 
* OUTPUT: fake_bl_108 
* OUTPUT: fake_br_108 
* OUTPUT: fake_bl_109 
* OUTPUT: fake_br_109 
* OUTPUT: fake_bl_110 
* OUTPUT: fake_br_110 
* OUTPUT: fake_bl_111 
* OUTPUT: fake_br_111 
* OUTPUT: fake_bl_112 
* OUTPUT: fake_br_112 
* OUTPUT: fake_bl_113 
* OUTPUT: fake_br_113 
* OUTPUT: fake_bl_114 
* OUTPUT: fake_br_114 
* OUTPUT: fake_bl_115 
* OUTPUT: fake_br_115 
* OUTPUT: fake_bl_116 
* OUTPUT: fake_br_116 
* OUTPUT: fake_bl_117 
* OUTPUT: fake_br_117 
* OUTPUT: fake_bl_118 
* OUTPUT: fake_br_118 
* OUTPUT: fake_bl_119 
* OUTPUT: fake_br_119 
* OUTPUT: fake_bl_120 
* OUTPUT: fake_br_120 
* OUTPUT: fake_bl_121 
* OUTPUT: fake_br_121 
* OUTPUT: fake_bl_122 
* OUTPUT: fake_br_122 
* OUTPUT: fake_bl_123 
* OUTPUT: fake_br_123 
* OUTPUT: fake_bl_124 
* OUTPUT: fake_br_124 
* OUTPUT: fake_bl_125 
* OUTPUT: fake_br_125 
* OUTPUT: fake_bl_126 
* OUTPUT: fake_br_126 
* OUTPUT: fake_bl_127 
* OUTPUT: fake_br_127 
* OUTPUT: fake_bl_128 
* OUTPUT: fake_br_128 
* POWER : vdd 
* GROUND: gnd 
* BIAS  : gate 
Xrca_top_0
+ fake_bl_0 vdd gnd fake_br_0 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_1
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_2
+ fake_bl_1 vdd gnd fake_br_1 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_3
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_4
+ fake_bl_2 vdd gnd fake_br_2 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_5
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_6
+ fake_bl_3 vdd gnd fake_br_3 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_7
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_8
+ fake_bl_4 vdd gnd fake_br_4 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_9
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_10
+ fake_bl_5 vdd gnd fake_br_5 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_11
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_12
+ fake_bl_6 vdd gnd fake_br_6 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_13
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_14
+ fake_bl_7 vdd gnd fake_br_7 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_15
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_16
+ fake_bl_8 vdd gnd fake_br_8 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_17
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_18
+ fake_bl_9 vdd gnd fake_br_9 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_19
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_20
+ fake_bl_10 vdd gnd fake_br_10 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_21
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_22
+ fake_bl_11 vdd gnd fake_br_11 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_23
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_24
+ fake_bl_12 vdd gnd fake_br_12 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_25
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_26
+ fake_bl_13 vdd gnd fake_br_13 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_27
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_28
+ fake_bl_14 vdd gnd fake_br_14 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_29
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_30
+ fake_bl_15 vdd gnd fake_br_15 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_31
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_32
+ fake_bl_16 vdd gnd fake_br_16 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_33
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_34
+ fake_bl_17 vdd gnd fake_br_17 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_35
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_36
+ fake_bl_18 vdd gnd fake_br_18 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_37
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_38
+ fake_bl_19 vdd gnd fake_br_19 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_39
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_40
+ fake_bl_20 vdd gnd fake_br_20 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_41
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_42
+ fake_bl_21 vdd gnd fake_br_21 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_43
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_44
+ fake_bl_22 vdd gnd fake_br_22 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_45
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_46
+ fake_bl_23 vdd gnd fake_br_23 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_47
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_48
+ fake_bl_24 vdd gnd fake_br_24 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_49
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_50
+ fake_bl_25 vdd gnd fake_br_25 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_51
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_52
+ fake_bl_26 vdd gnd fake_br_26 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_53
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_54
+ fake_bl_27 vdd gnd fake_br_27 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_55
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_56
+ fake_bl_28 vdd gnd fake_br_28 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_57
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_58
+ fake_bl_29 vdd gnd fake_br_29 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_59
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_60
+ fake_bl_30 vdd gnd fake_br_30 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_61
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_62
+ fake_bl_31 vdd gnd fake_br_31 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_63
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_64
+ fake_bl_32 vdd gnd fake_br_32 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_65
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_66
+ fake_bl_33 vdd gnd fake_br_33 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_67
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_68
+ fake_bl_34 vdd gnd fake_br_34 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_69
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_70
+ fake_bl_35 vdd gnd fake_br_35 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_71
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_72
+ fake_bl_36 vdd gnd fake_br_36 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_73
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_74
+ fake_bl_37 vdd gnd fake_br_37 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_75
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_76
+ fake_bl_38 vdd gnd fake_br_38 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_77
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_78
+ fake_bl_39 vdd gnd fake_br_39 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_79
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_80
+ fake_bl_40 vdd gnd fake_br_40 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_81
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_82
+ fake_bl_41 vdd gnd fake_br_41 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_83
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_84
+ fake_bl_42 vdd gnd fake_br_42 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_85
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_86
+ fake_bl_43 vdd gnd fake_br_43 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_87
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_88
+ fake_bl_44 vdd gnd fake_br_44 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_89
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_90
+ fake_bl_45 vdd gnd fake_br_45 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_91
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_92
+ fake_bl_46 vdd gnd fake_br_46 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_93
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_94
+ fake_bl_47 vdd gnd fake_br_47 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_95
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_96
+ fake_bl_48 vdd gnd fake_br_48 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_97
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_98
+ fake_bl_49 vdd gnd fake_br_49 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_99
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_100
+ fake_bl_50 vdd gnd fake_br_50 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_101
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_102
+ fake_bl_51 vdd gnd fake_br_51 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_103
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_104
+ fake_bl_52 vdd gnd fake_br_52 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_105
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_106
+ fake_bl_53 vdd gnd fake_br_53 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_107
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_108
+ fake_bl_54 vdd gnd fake_br_54 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_109
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_110
+ fake_bl_55 vdd gnd fake_br_55 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_111
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_112
+ fake_bl_56 vdd gnd fake_br_56 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_113
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_114
+ fake_bl_57 vdd gnd fake_br_57 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_115
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_116
+ fake_bl_58 vdd gnd fake_br_58 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_117
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_118
+ fake_bl_59 vdd gnd fake_br_59 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_119
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_120
+ fake_bl_60 vdd gnd fake_br_60 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_121
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_122
+ fake_bl_61 vdd gnd fake_br_61 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_123
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_124
+ fake_bl_62 vdd gnd fake_br_62 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_125
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_126
+ fake_bl_63 vdd gnd fake_br_63 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_127
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_128
+ fake_bl_64 vdd gnd fake_br_64 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_129
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_130
+ fake_bl_65 vdd gnd fake_br_65 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_131
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_132
+ fake_bl_66 vdd gnd fake_br_66 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_133
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_134
+ fake_bl_67 vdd gnd fake_br_67 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_135
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_136
+ fake_bl_68 vdd gnd fake_br_68 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_137
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_138
+ fake_bl_69 vdd gnd fake_br_69 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_139
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_140
+ fake_bl_70 vdd gnd fake_br_70 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_141
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_142
+ fake_bl_71 vdd gnd fake_br_71 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_143
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_144
+ fake_bl_72 vdd gnd fake_br_72 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_145
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_146
+ fake_bl_73 vdd gnd fake_br_73 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_147
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_148
+ fake_bl_74 vdd gnd fake_br_74 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_149
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_150
+ fake_bl_75 vdd gnd fake_br_75 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_151
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_152
+ fake_bl_76 vdd gnd fake_br_76 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_153
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_154
+ fake_bl_77 vdd gnd fake_br_77 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_155
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_156
+ fake_bl_78 vdd gnd fake_br_78 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_157
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_158
+ fake_bl_79 vdd gnd fake_br_79 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_159
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_160
+ fake_bl_80 vdd gnd fake_br_80 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_161
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_162
+ fake_bl_81 vdd gnd fake_br_81 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_163
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_164
+ fake_bl_82 vdd gnd fake_br_82 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_165
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_166
+ fake_bl_83 vdd gnd fake_br_83 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_167
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_168
+ fake_bl_84 vdd gnd fake_br_84 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_169
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_170
+ fake_bl_85 vdd gnd fake_br_85 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_171
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_172
+ fake_bl_86 vdd gnd fake_br_86 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_173
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_174
+ fake_bl_87 vdd gnd fake_br_87 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_175
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_176
+ fake_bl_88 vdd gnd fake_br_88 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_177
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_178
+ fake_bl_89 vdd gnd fake_br_89 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_179
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_180
+ fake_bl_90 vdd gnd fake_br_90 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_181
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_182
+ fake_bl_91 vdd gnd fake_br_91 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_183
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_184
+ fake_bl_92 vdd gnd fake_br_92 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_185
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_186
+ fake_bl_93 vdd gnd fake_br_93 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_187
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_188
+ fake_bl_94 vdd gnd fake_br_94 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_189
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_190
+ fake_bl_95 vdd gnd fake_br_95 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_191
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_192
+ fake_bl_96 vdd gnd fake_br_96 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_193
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_194
+ fake_bl_97 vdd gnd fake_br_97 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_195
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_196
+ fake_bl_98 vdd gnd fake_br_98 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_197
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_198
+ fake_bl_99 vdd gnd fake_br_99 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_199
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_200
+ fake_bl_100 vdd gnd fake_br_100 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_201
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_202
+ fake_bl_101 vdd gnd fake_br_101 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_203
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_204
+ fake_bl_102 vdd gnd fake_br_102 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_205
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_206
+ fake_bl_103 vdd gnd fake_br_103 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_207
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_208
+ fake_bl_104 vdd gnd fake_br_104 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_209
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_210
+ fake_bl_105 vdd gnd fake_br_105 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_211
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_212
+ fake_bl_106 vdd gnd fake_br_106 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_213
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_214
+ fake_bl_107 vdd gnd fake_br_107 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_215
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_216
+ fake_bl_108 vdd gnd fake_br_108 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_217
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_218
+ fake_bl_109 vdd gnd fake_br_109 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_219
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_220
+ fake_bl_110 vdd gnd fake_br_110 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_221
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_222
+ fake_bl_111 vdd gnd fake_br_111 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_223
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_224
+ fake_bl_112 vdd gnd fake_br_112 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_225
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_226
+ fake_bl_113 vdd gnd fake_br_113 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_227
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_228
+ fake_bl_114 vdd gnd fake_br_114 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_229
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_230
+ fake_bl_115 vdd gnd fake_br_115 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_231
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_232
+ fake_bl_116 vdd gnd fake_br_116 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_233
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_234
+ fake_bl_117 vdd gnd fake_br_117 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_235
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_236
+ fake_bl_118 vdd gnd fake_br_118 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_237
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_238
+ fake_bl_119 vdd gnd fake_br_119 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_239
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_240
+ fake_bl_120 vdd gnd fake_br_120 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_241
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_242
+ fake_bl_121 vdd gnd fake_br_121 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_243
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_244
+ fake_bl_122 vdd gnd fake_br_122 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_245
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_246
+ fake_bl_123 vdd gnd fake_br_123 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_247
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_248
+ fake_bl_124 vdd gnd fake_br_124 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_249
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_250
+ fake_bl_125 vdd gnd fake_br_125 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_251
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_252
+ fake_bl_126 vdd gnd fake_br_126 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_253
+ vdd vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend_cent
Xrca_top_254
+ fake_bl_127 vdd gnd fake_br_127 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
Xrca_top_255
+ gnd vdd vnb
+ sky130_fd_bd_sram__sram_sp_colend_p_cent
Xrca_top_256
+ fake_bl_128 vdd gnd fake_br_128 gate vdd gnd
+ sky130_fd_bd_sram__sram_sp_colend
.ENDS sky130_sram_1kbyte_1rw_32x256_8_sky130_col_cap_array
* NGSPICE file created from sky130_fd_bd_sram__openram_sp_rowend_replica.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_rowend_replica VPWR WL
.ends
* NGSPICE file created from sky130_fd_bd_sram__sram_sp_corner.ext - technology: sky130A

.subckt sky130_fd_bd_sram__sram_sp_corner VPWR VPB VNB
.ends
* NGSPICE file created from sky130_fd_bd_sram__openram_sp_rowenda_replica.ext - technology: sky130A

.subckt sky130_fd_bd_sram__openram_sp_rowenda_replica VPWR WL
.ends

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_sky130_row_cap_array
+ wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9
+ wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17
+ wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25
+ wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33
+ wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41
+ wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49
+ wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57
+ wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 wl_0_65
+ wl_0_66 wl_0_67 vdd gnd
* OUTPUT: wl_0_0 
* OUTPUT: wl_0_1 
* OUTPUT: wl_0_2 
* OUTPUT: wl_0_3 
* OUTPUT: wl_0_4 
* OUTPUT: wl_0_5 
* OUTPUT: wl_0_6 
* OUTPUT: wl_0_7 
* OUTPUT: wl_0_8 
* OUTPUT: wl_0_9 
* OUTPUT: wl_0_10 
* OUTPUT: wl_0_11 
* OUTPUT: wl_0_12 
* OUTPUT: wl_0_13 
* OUTPUT: wl_0_14 
* OUTPUT: wl_0_15 
* OUTPUT: wl_0_16 
* OUTPUT: wl_0_17 
* OUTPUT: wl_0_18 
* OUTPUT: wl_0_19 
* OUTPUT: wl_0_20 
* OUTPUT: wl_0_21 
* OUTPUT: wl_0_22 
* OUTPUT: wl_0_23 
* OUTPUT: wl_0_24 
* OUTPUT: wl_0_25 
* OUTPUT: wl_0_26 
* OUTPUT: wl_0_27 
* OUTPUT: wl_0_28 
* OUTPUT: wl_0_29 
* OUTPUT: wl_0_30 
* OUTPUT: wl_0_31 
* OUTPUT: wl_0_32 
* OUTPUT: wl_0_33 
* OUTPUT: wl_0_34 
* OUTPUT: wl_0_35 
* OUTPUT: wl_0_36 
* OUTPUT: wl_0_37 
* OUTPUT: wl_0_38 
* OUTPUT: wl_0_39 
* OUTPUT: wl_0_40 
* OUTPUT: wl_0_41 
* OUTPUT: wl_0_42 
* OUTPUT: wl_0_43 
* OUTPUT: wl_0_44 
* OUTPUT: wl_0_45 
* OUTPUT: wl_0_46 
* OUTPUT: wl_0_47 
* OUTPUT: wl_0_48 
* OUTPUT: wl_0_49 
* OUTPUT: wl_0_50 
* OUTPUT: wl_0_51 
* OUTPUT: wl_0_52 
* OUTPUT: wl_0_53 
* OUTPUT: wl_0_54 
* OUTPUT: wl_0_55 
* OUTPUT: wl_0_56 
* OUTPUT: wl_0_57 
* OUTPUT: wl_0_58 
* OUTPUT: wl_0_59 
* OUTPUT: wl_0_60 
* OUTPUT: wl_0_61 
* OUTPUT: wl_0_62 
* OUTPUT: wl_0_63 
* OUTPUT: wl_0_64 
* OUTPUT: wl_0_65 
* OUTPUT: wl_0_66 
* OUTPUT: wl_0_67 
* POWER : vdd 
* GROUND: gnd 
Xrca_0
+ vdd gnd vdd
+ sky130_fd_bd_sram__sram_sp_cornera
Xrca_1
+ wl_0_0 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_2
+ wl_0_1 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_3
+ wl_0_2 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_4
+ wl_0_3 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_5
+ wl_0_4 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_6
+ wl_0_5 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_7
+ wl_0_6 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_8
+ wl_0_7 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_9
+ wl_0_8 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_10
+ wl_0_9 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_11
+ wl_0_10 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_12
+ wl_0_11 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_13
+ wl_0_12 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_14
+ wl_0_13 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_15
+ wl_0_14 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_16
+ wl_0_15 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_17
+ wl_0_16 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_18
+ wl_0_17 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_19
+ wl_0_18 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_20
+ wl_0_19 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_21
+ wl_0_20 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_22
+ wl_0_21 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_23
+ wl_0_22 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_24
+ wl_0_23 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_25
+ wl_0_24 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_26
+ wl_0_25 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_27
+ wl_0_26 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_28
+ wl_0_27 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_29
+ wl_0_28 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_30
+ wl_0_29 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_31
+ wl_0_30 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_32
+ wl_0_31 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_33
+ wl_0_32 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_34
+ wl_0_33 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_35
+ wl_0_34 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_36
+ wl_0_35 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_37
+ wl_0_36 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_38
+ wl_0_37 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_39
+ wl_0_38 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_40
+ wl_0_39 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_41
+ wl_0_40 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_42
+ wl_0_41 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_43
+ wl_0_42 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_44
+ wl_0_43 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_45
+ wl_0_44 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_46
+ wl_0_45 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_47
+ wl_0_46 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_48
+ wl_0_47 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_49
+ wl_0_48 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_50
+ wl_0_49 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_51
+ wl_0_50 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_52
+ wl_0_51 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_53
+ wl_0_52 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_54
+ wl_0_53 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_55
+ wl_0_54 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_56
+ wl_0_55 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_57
+ wl_0_56 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_58
+ wl_0_57 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_59
+ wl_0_58 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_60
+ wl_0_59 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_61
+ wl_0_60 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_62
+ wl_0_61 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_63
+ wl_0_62 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_64
+ wl_0_63 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_65
+ wl_0_64 vdd
+ sky130_fd_bd_sram__openram_sp_rowenda_replica
Xrca_66
+ wl_0_65 vdd
+ sky130_fd_bd_sram__openram_sp_rowend_replica
Xrca_67
+ vdd gnd vdd
+ sky130_fd_bd_sram__sram_sp_corner
.ENDS sky130_sram_1kbyte_1rw_32x256_8_sky130_row_cap_array

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_sky130_replica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48
+ wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56
+ wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 vdd
+ gnd
* INOUT : rbl_bl_0_0 
* INOUT : rbl_br_0_0 
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INPUT : rbl_wl_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* POWER : vdd 
* GROUND: gnd 
* rows: 65 cols: 129
* rbl: [1, 0] left_rbl: [0] right_rbl: []
Xbitcell_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 wl_0_0 wl_0_1 wl_0_2
+ wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11
+ wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19
+ wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27
+ wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35
+ wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43
+ wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51
+ wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59
+ wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_sky130_bitcell_array
Xreplica_col_0
+ rbl_bl_0_0 rbl_br_0_0 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4
+ wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13
+ wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21
+ wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29
+ wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37
+ wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45
+ wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53
+ wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61
+ wl_0_62 wl_0_63 wl_0_64 vdd gnd gnd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_sky130_replica_column
Xdummy_row_0
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 rbl_wl_0_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_sky130_dummy_array
Xdummy_row_bot
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 vdd gnd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_sky130_col_cap_array_0
Xdummy_row_top
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 bl_0_65 br_0_65
+ bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68 bl_0_69 br_0_69
+ bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72 bl_0_73 br_0_73
+ bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76 bl_0_77 br_0_77
+ bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80 bl_0_81 br_0_81
+ bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84 bl_0_85 br_0_85
+ bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88 bl_0_89 br_0_89
+ bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92 bl_0_93 br_0_93
+ bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96 bl_0_97 br_0_97
+ bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100 bl_0_101 br_0_101
+ bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104 br_0_104 bl_0_105
+ br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107 bl_0_108 br_0_108
+ bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111 br_0_111 bl_0_112
+ br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114 bl_0_115 br_0_115
+ bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118 br_0_118 bl_0_119
+ br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121 bl_0_122 br_0_122
+ bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125 br_0_125 bl_0_126
+ br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 vdd gnd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_sky130_col_cap_array
Xdummy_col_left
+ gnd rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48
+ wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56
+ wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 gnd
+ vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_sky130_row_cap_array
Xdummy_col_right
+ gnd rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48
+ wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56
+ wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 gnd
+ vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_sky130_row_cap_array_0
.ENDS sky130_sram_1kbyte_1rw_32x256_8_sky130_replica_bitcell_array

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_sky130_capped_replica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48
+ wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56
+ wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 vdd
+ gnd
* INOUT : rbl_bl_0_0 
* INOUT : rbl_br_0_0 
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INOUT : bl_0_65 
* INOUT : br_0_65 
* INOUT : bl_0_66 
* INOUT : br_0_66 
* INOUT : bl_0_67 
* INOUT : br_0_67 
* INOUT : bl_0_68 
* INOUT : br_0_68 
* INOUT : bl_0_69 
* INOUT : br_0_69 
* INOUT : bl_0_70 
* INOUT : br_0_70 
* INOUT : bl_0_71 
* INOUT : br_0_71 
* INOUT : bl_0_72 
* INOUT : br_0_72 
* INOUT : bl_0_73 
* INOUT : br_0_73 
* INOUT : bl_0_74 
* INOUT : br_0_74 
* INOUT : bl_0_75 
* INOUT : br_0_75 
* INOUT : bl_0_76 
* INOUT : br_0_76 
* INOUT : bl_0_77 
* INOUT : br_0_77 
* INOUT : bl_0_78 
* INOUT : br_0_78 
* INOUT : bl_0_79 
* INOUT : br_0_79 
* INOUT : bl_0_80 
* INOUT : br_0_80 
* INOUT : bl_0_81 
* INOUT : br_0_81 
* INOUT : bl_0_82 
* INOUT : br_0_82 
* INOUT : bl_0_83 
* INOUT : br_0_83 
* INOUT : bl_0_84 
* INOUT : br_0_84 
* INOUT : bl_0_85 
* INOUT : br_0_85 
* INOUT : bl_0_86 
* INOUT : br_0_86 
* INOUT : bl_0_87 
* INOUT : br_0_87 
* INOUT : bl_0_88 
* INOUT : br_0_88 
* INOUT : bl_0_89 
* INOUT : br_0_89 
* INOUT : bl_0_90 
* INOUT : br_0_90 
* INOUT : bl_0_91 
* INOUT : br_0_91 
* INOUT : bl_0_92 
* INOUT : br_0_92 
* INOUT : bl_0_93 
* INOUT : br_0_93 
* INOUT : bl_0_94 
* INOUT : br_0_94 
* INOUT : bl_0_95 
* INOUT : br_0_95 
* INOUT : bl_0_96 
* INOUT : br_0_96 
* INOUT : bl_0_97 
* INOUT : br_0_97 
* INOUT : bl_0_98 
* INOUT : br_0_98 
* INOUT : bl_0_99 
* INOUT : br_0_99 
* INOUT : bl_0_100 
* INOUT : br_0_100 
* INOUT : bl_0_101 
* INOUT : br_0_101 
* INOUT : bl_0_102 
* INOUT : br_0_102 
* INOUT : bl_0_103 
* INOUT : br_0_103 
* INOUT : bl_0_104 
* INOUT : br_0_104 
* INOUT : bl_0_105 
* INOUT : br_0_105 
* INOUT : bl_0_106 
* INOUT : br_0_106 
* INOUT : bl_0_107 
* INOUT : br_0_107 
* INOUT : bl_0_108 
* INOUT : br_0_108 
* INOUT : bl_0_109 
* INOUT : br_0_109 
* INOUT : bl_0_110 
* INOUT : br_0_110 
* INOUT : bl_0_111 
* INOUT : br_0_111 
* INOUT : bl_0_112 
* INOUT : br_0_112 
* INOUT : bl_0_113 
* INOUT : br_0_113 
* INOUT : bl_0_114 
* INOUT : br_0_114 
* INOUT : bl_0_115 
* INOUT : br_0_115 
* INOUT : bl_0_116 
* INOUT : br_0_116 
* INOUT : bl_0_117 
* INOUT : br_0_117 
* INOUT : bl_0_118 
* INOUT : br_0_118 
* INOUT : bl_0_119 
* INOUT : br_0_119 
* INOUT : bl_0_120 
* INOUT : br_0_120 
* INOUT : bl_0_121 
* INOUT : br_0_121 
* INOUT : bl_0_122 
* INOUT : br_0_122 
* INOUT : bl_0_123 
* INOUT : br_0_123 
* INOUT : bl_0_124 
* INOUT : br_0_124 
* INOUT : bl_0_125 
* INOUT : br_0_125 
* INOUT : bl_0_126 
* INOUT : br_0_126 
* INOUT : bl_0_127 
* INOUT : br_0_127 
* INOUT : bl_0_128 
* INOUT : br_0_128 
* INPUT : rbl_wl_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* POWER : vdd 
* GROUND: gnd 
* rows: 65 cols: 129
* rbl: [1, 0] left_rbl: [0] right_rbl: []
Xreplica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128
+ rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48
+ wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56
+ wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 vdd
+ gnd
+ sky130_sram_1kbyte_1rw_32x256_8_sky130_replica_bitcell_array
.ENDS sky130_sram_1kbyte_1rw_32x256_8_sky130_capped_replica_bitcell_array

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_bank
+ dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7
+ dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15
+ dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22
+ dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29
+ dout0_30 dout0_31 dout0_32 rbl_bl_0_0 din0_0 din0_1 din0_2 din0_3
+ din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12
+ din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20
+ din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28
+ din0_29 din0_30 din0_31 din0_32 addr0_0 addr0_1 addr0_2 addr0_3
+ addr0_4 addr0_5 addr0_6 addr0_7 addr0_8 s_en0 p_en_bar0 w_en0
+ bank_wmask0_0 bank_wmask0_1 bank_wmask0_2 bank_wmask0_3
+ bank_spare_wen0_0 wl_en0 vdd gnd
* OUTPUT: dout0_0 
* OUTPUT: dout0_1 
* OUTPUT: dout0_2 
* OUTPUT: dout0_3 
* OUTPUT: dout0_4 
* OUTPUT: dout0_5 
* OUTPUT: dout0_6 
* OUTPUT: dout0_7 
* OUTPUT: dout0_8 
* OUTPUT: dout0_9 
* OUTPUT: dout0_10 
* OUTPUT: dout0_11 
* OUTPUT: dout0_12 
* OUTPUT: dout0_13 
* OUTPUT: dout0_14 
* OUTPUT: dout0_15 
* OUTPUT: dout0_16 
* OUTPUT: dout0_17 
* OUTPUT: dout0_18 
* OUTPUT: dout0_19 
* OUTPUT: dout0_20 
* OUTPUT: dout0_21 
* OUTPUT: dout0_22 
* OUTPUT: dout0_23 
* OUTPUT: dout0_24 
* OUTPUT: dout0_25 
* OUTPUT: dout0_26 
* OUTPUT: dout0_27 
* OUTPUT: dout0_28 
* OUTPUT: dout0_29 
* OUTPUT: dout0_30 
* OUTPUT: dout0_31 
* OUTPUT: dout0_32 
* OUTPUT: rbl_bl_0_0 
* INPUT : din0_0 
* INPUT : din0_1 
* INPUT : din0_2 
* INPUT : din0_3 
* INPUT : din0_4 
* INPUT : din0_5 
* INPUT : din0_6 
* INPUT : din0_7 
* INPUT : din0_8 
* INPUT : din0_9 
* INPUT : din0_10 
* INPUT : din0_11 
* INPUT : din0_12 
* INPUT : din0_13 
* INPUT : din0_14 
* INPUT : din0_15 
* INPUT : din0_16 
* INPUT : din0_17 
* INPUT : din0_18 
* INPUT : din0_19 
* INPUT : din0_20 
* INPUT : din0_21 
* INPUT : din0_22 
* INPUT : din0_23 
* INPUT : din0_24 
* INPUT : din0_25 
* INPUT : din0_26 
* INPUT : din0_27 
* INPUT : din0_28 
* INPUT : din0_29 
* INPUT : din0_30 
* INPUT : din0_31 
* INPUT : din0_32 
* INPUT : addr0_0 
* INPUT : addr0_1 
* INPUT : addr0_2 
* INPUT : addr0_3 
* INPUT : addr0_4 
* INPUT : addr0_5 
* INPUT : addr0_6 
* INPUT : addr0_7 
* INPUT : addr0_8 
* INPUT : s_en0 
* INPUT : p_en_bar0 
* INPUT : w_en0 
* INPUT : bank_wmask0_0 
* INPUT : bank_wmask0_1 
* INPUT : bank_wmask0_2 
* INPUT : bank_wmask0_3 
* INPUT : bank_spare_wen0_0 
* INPUT : wl_en0 
* POWER : vdd 
* GROUND: gnd 
Xbitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 rbl_wl0
+ wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9
+ wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17
+ wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25
+ wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33
+ wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41
+ wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49
+ wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57
+ wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_sky130_capped_replica_bitcell_array
Xport_data0
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64
+ bl_0_65 br_0_65 bl_0_66 br_0_66 bl_0_67 br_0_67 bl_0_68 br_0_68
+ bl_0_69 br_0_69 bl_0_70 br_0_70 bl_0_71 br_0_71 bl_0_72 br_0_72
+ bl_0_73 br_0_73 bl_0_74 br_0_74 bl_0_75 br_0_75 bl_0_76 br_0_76
+ bl_0_77 br_0_77 bl_0_78 br_0_78 bl_0_79 br_0_79 bl_0_80 br_0_80
+ bl_0_81 br_0_81 bl_0_82 br_0_82 bl_0_83 br_0_83 bl_0_84 br_0_84
+ bl_0_85 br_0_85 bl_0_86 br_0_86 bl_0_87 br_0_87 bl_0_88 br_0_88
+ bl_0_89 br_0_89 bl_0_90 br_0_90 bl_0_91 br_0_91 bl_0_92 br_0_92
+ bl_0_93 br_0_93 bl_0_94 br_0_94 bl_0_95 br_0_95 bl_0_96 br_0_96
+ bl_0_97 br_0_97 bl_0_98 br_0_98 bl_0_99 br_0_99 bl_0_100 br_0_100
+ bl_0_101 br_0_101 bl_0_102 br_0_102 bl_0_103 br_0_103 bl_0_104
+ br_0_104 bl_0_105 br_0_105 bl_0_106 br_0_106 bl_0_107 br_0_107
+ bl_0_108 br_0_108 bl_0_109 br_0_109 bl_0_110 br_0_110 bl_0_111
+ br_0_111 bl_0_112 br_0_112 bl_0_113 br_0_113 bl_0_114 br_0_114
+ bl_0_115 br_0_115 bl_0_116 br_0_116 bl_0_117 br_0_117 bl_0_118
+ br_0_118 bl_0_119 br_0_119 bl_0_120 br_0_120 bl_0_121 br_0_121
+ bl_0_122 br_0_122 bl_0_123 br_0_123 bl_0_124 br_0_124 bl_0_125
+ br_0_125 bl_0_126 br_0_126 bl_0_127 br_0_127 bl_0_128 br_0_128 dout0_0
+ dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8
+ dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16
+ dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23
+ dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30
+ dout0_31 dout0_32 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6
+ din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15
+ din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23
+ din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31
+ din0_32 sel0_0 sel0_1 sel0_2 sel0_3 s_en0 p_en_bar0 w_en0
+ bank_wmask0_0 bank_wmask0_1 bank_wmask0_2 bank_wmask0_3
+ bank_spare_wen0_0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_port_data
Xport_address0
+ addr0_2 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 addr0_8 wl_en0 wl_0_0
+ wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 wl_0_33 wl_0_34
+ wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40 wl_0_41 wl_0_42
+ wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48 wl_0_49 wl_0_50
+ wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56 wl_0_57 wl_0_58
+ wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64 rbl_wl0 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_port_address
Xcol_address_decoder0
+ addr0_0 addr0_1 sel0_0 sel0_1 sel0_2 sel0_3 vdd gnd
+ sky130_sram_1kbyte_1rw_32x256_8_column_decoder
.ENDS sky130_sram_1kbyte_1rw_32x256_8_bank

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_row_addr_dff
+ din_0 din_1 din_2 din_3 din_4 din_5 din_6 dout_0 dout_1 dout_2 dout_3
+ dout_4 dout_5 dout_6 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 7 cols: 1
Xdff_r0_c0
+ din_0 dout_0 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r1_c0
+ din_1 dout_1 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r2_c0
+ din_2 dout_2 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r3_c0
+ din_3 dout_3 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r4_c0
+ din_4 dout_4 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r5_c0
+ din_5 dout_5 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r6_c0
+ din_6 dout_6 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
.ENDS sky130_sram_1kbyte_1rw_32x256_8_row_addr_dff

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8_data_dff
+ din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10
+ din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20
+ din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30
+ din_31 din_32 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7
+ dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16
+ dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24
+ dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 dout_32 clk
+ vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : din_32 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* OUTPUT: dout_32 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 33
Xdff_r0_c0
+ din_0 dout_0 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c1
+ din_1 dout_1 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c2
+ din_2 dout_2 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c3
+ din_3 dout_3 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c4
+ din_4 dout_4 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c5
+ din_5 dout_5 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c6
+ din_6 dout_6 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c7
+ din_7 dout_7 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c8
+ din_8 dout_8 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c9
+ din_9 dout_9 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c10
+ din_10 dout_10 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c11
+ din_11 dout_11 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c12
+ din_12 dout_12 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c13
+ din_13 dout_13 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c14
+ din_14 dout_14 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c15
+ din_15 dout_15 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c16
+ din_16 dout_16 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c17
+ din_17 dout_17 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c18
+ din_18 dout_18 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c19
+ din_19 dout_19 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c20
+ din_20 dout_20 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c21
+ din_21 dout_21 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c22
+ din_22 dout_22 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c23
+ din_23 dout_23 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c24
+ din_24 dout_24 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c25
+ din_25 dout_25 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c26
+ din_26 dout_26 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c27
+ din_27 dout_27 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c28
+ din_28 dout_28 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c29
+ din_29 dout_29 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c30
+ din_30 dout_30 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c31
+ din_31 dout_31 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
Xdff_r0_c32
+ din_32 dout_32 CLK VDD GND
+ sky130_fd_bd_sram__openram_dff
.ENDS sky130_sram_1kbyte_1rw_32x256_8_data_dff

.SUBCKT sky130_sram_1kbyte_1rw_32x256_8
+ din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7]
+ din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22]
+ din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29]
+ din0[30] din0[31] din0[32] addr0[0] addr0[1] addr0[2] addr0[3]
+ addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] csb0 web0 clk0 wmask0[0]
+ wmask0[1] wmask0[2] wmask0[3] spare_wen0 dout0[0] dout0[1] dout0[2]
+ dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9]
+ dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16]
+ dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23]
+ dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30]
+ dout0[31] dout0[32] vccd1 vssd1
* INPUT : din0[0] 
* INPUT : din0[1] 
* INPUT : din0[2] 
* INPUT : din0[3] 
* INPUT : din0[4] 
* INPUT : din0[5] 
* INPUT : din0[6] 
* INPUT : din0[7] 
* INPUT : din0[8] 
* INPUT : din0[9] 
* INPUT : din0[10] 
* INPUT : din0[11] 
* INPUT : din0[12] 
* INPUT : din0[13] 
* INPUT : din0[14] 
* INPUT : din0[15] 
* INPUT : din0[16] 
* INPUT : din0[17] 
* INPUT : din0[18] 
* INPUT : din0[19] 
* INPUT : din0[20] 
* INPUT : din0[21] 
* INPUT : din0[22] 
* INPUT : din0[23] 
* INPUT : din0[24] 
* INPUT : din0[25] 
* INPUT : din0[26] 
* INPUT : din0[27] 
* INPUT : din0[28] 
* INPUT : din0[29] 
* INPUT : din0[30] 
* INPUT : din0[31] 
* INPUT : din0[32] 
* INPUT : addr0[0] 
* INPUT : addr0[1] 
* INPUT : addr0[2] 
* INPUT : addr0[3] 
* INPUT : addr0[4] 
* INPUT : addr0[5] 
* INPUT : addr0[6] 
* INPUT : addr0[7] 
* INPUT : addr0[8] 
* INPUT : csb0 
* INPUT : web0 
* INPUT : clk0 
* INPUT : wmask0[0] 
* INPUT : wmask0[1] 
* INPUT : wmask0[2] 
* INPUT : wmask0[3] 
* INPUT : spare_wen0 
* OUTPUT: dout0[0] 
* OUTPUT: dout0[1] 
* OUTPUT: dout0[2] 
* OUTPUT: dout0[3] 
* OUTPUT: dout0[4] 
* OUTPUT: dout0[5] 
* OUTPUT: dout0[6] 
* OUTPUT: dout0[7] 
* OUTPUT: dout0[8] 
* OUTPUT: dout0[9] 
* OUTPUT: dout0[10] 
* OUTPUT: dout0[11] 
* OUTPUT: dout0[12] 
* OUTPUT: dout0[13] 
* OUTPUT: dout0[14] 
* OUTPUT: dout0[15] 
* OUTPUT: dout0[16] 
* OUTPUT: dout0[17] 
* OUTPUT: dout0[18] 
* OUTPUT: dout0[19] 
* OUTPUT: dout0[20] 
* OUTPUT: dout0[21] 
* OUTPUT: dout0[22] 
* OUTPUT: dout0[23] 
* OUTPUT: dout0[24] 
* OUTPUT: dout0[25] 
* OUTPUT: dout0[26] 
* OUTPUT: dout0[27] 
* OUTPUT: dout0[28] 
* OUTPUT: dout0[29] 
* OUTPUT: dout0[30] 
* OUTPUT: dout0[31] 
* OUTPUT: dout0[32] 
* POWER : vccd1 
* GROUND: vssd1 
Xbank0
+ dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6]
+ dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13]
+ dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20]
+ dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[30] dout0[31] dout0[32] rbl_bl0 bank_din0_0
+ bank_din0_1 bank_din0_2 bank_din0_3 bank_din0_4 bank_din0_5
+ bank_din0_6 bank_din0_7 bank_din0_8 bank_din0_9 bank_din0_10
+ bank_din0_11 bank_din0_12 bank_din0_13 bank_din0_14 bank_din0_15
+ bank_din0_16 bank_din0_17 bank_din0_18 bank_din0_19 bank_din0_20
+ bank_din0_21 bank_din0_22 bank_din0_23 bank_din0_24 bank_din0_25
+ bank_din0_26 bank_din0_27 bank_din0_28 bank_din0_29 bank_din0_30
+ bank_din0_31 bank_din0_32 a0_0 a0_1 a0_2 a0_3 a0_4 a0_5 a0_6 a0_7 a0_8
+ s_en0 p_en_bar0 w_en0 bank_wmask0_0 bank_wmask0_1 bank_wmask0_2
+ bank_wmask0_3 bank_spare_wen0_0 wl_en0 vccd1 vssd1
+ sky130_sram_1kbyte_1rw_32x256_8_bank
Xcontrol0
+ csb0 web0 clk0 rbl_bl0 s_en0 w_en0 p_en_bar0 wl_en0 clk_buf0 vccd1
+ vssd1
+ sky130_sram_1kbyte_1rw_32x256_8_control_logic_rw
Xrow_address0
+ addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] a0_2
+ a0_3 a0_4 a0_5 a0_6 a0_7 a0_8 clk_buf0 vccd1 vssd1
+ sky130_sram_1kbyte_1rw_32x256_8_row_addr_dff
Xcol_address0
+ addr0[0] addr0[1] a0_0 a0_1 clk_buf0 vccd1 vssd1
+ sky130_sram_1kbyte_1rw_32x256_8_col_addr_dff
Xwmask_dff0
+ wmask0[0] wmask0[1] wmask0[2] wmask0[3] bank_wmask0_0 bank_wmask0_1
+ bank_wmask0_2 bank_wmask0_3 clk_buf0 vccd1 vssd1
+ sky130_sram_1kbyte_1rw_32x256_8_wmask_dff
Xdata_dff0
+ din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7]
+ din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22]
+ din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29]
+ din0[30] din0[31] din0[32] bank_din0_0 bank_din0_1 bank_din0_2
+ bank_din0_3 bank_din0_4 bank_din0_5 bank_din0_6 bank_din0_7
+ bank_din0_8 bank_din0_9 bank_din0_10 bank_din0_11 bank_din0_12
+ bank_din0_13 bank_din0_14 bank_din0_15 bank_din0_16 bank_din0_17
+ bank_din0_18 bank_din0_19 bank_din0_20 bank_din0_21 bank_din0_22
+ bank_din0_23 bank_din0_24 bank_din0_25 bank_din0_26 bank_din0_27
+ bank_din0_28 bank_din0_29 bank_din0_30 bank_din0_31 bank_din0_32
+ clk_buf0 vccd1 vssd1
+ sky130_sram_1kbyte_1rw_32x256_8_data_dff
Xspare_wen_dff0
+ spare_wen0[0] bank_spare_wen0_0 clk_buf0 vccd1 vssd1
+ sky130_sram_1kbyte_1rw_32x256_8_spare_wen_dff
.ENDS sky130_sram_1kbyte_1rw_32x256_8
